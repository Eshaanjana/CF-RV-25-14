Stage5.bsv
// See LICENSE.iitm for license details
/*
Author: IIT Madras
Created on: Monday 21 June 2021 09:07:59 PM

*/
/*doc:overview:
This is the write-back stage of the pipeline where all instructions retire. By the time an
instructino reaches this stage it has been narrowed down via some of the previous stages into one of
the following categories of operations that can be performed in this stage:

  - SYSTEM: either xRET operations or CSR access operations.
  - TRAP: The instruction has encountered a trap during its operation in one of the previous stages.
  - BASEOUT: The instruction retirement includes a simple update to the registerfile
  - MEMOP: The instruction is either a cached store/atomic operation or an non-cached/IO memory op.

Each of the above have a unique ISB feeding in respective instructions to this module. This module
uses the fuid from the previous stage,  which maintains the order of instructions to find out which
ISB must be polled for the retiring/committing the next instruction.

Operations which can take multiple cycles in this stage are : CSR operations if daisy-chain is more
than 1 level deep; IO/non-cached Memory Operations may also take significantly longer in this stage
to complete.

All other ops will take a single cycle to complete.

When in simulation mode, this module will offload the commit-log packet to the test-bench via a
single Default-Reg (DReg) interface.

This module also instantiates the csrbox module, which hosts all the csrs and also the routines to
perform a trap or an xRet operation. Certain csr interfaces are simply bypassed along this module so
that they are exposed at the next hiegher level to rest of the pipeline and design.

*/
package stage5 ;

import FIFOF        :: * ;
import Vector       :: * ;
`ifdef async_rst
import SpecialFIFOs_Modified :: * ;
`else
import SpecialFIFOs :: * ;
`endif
import FIFOF        :: * ;
import TxRx         :: * ;
import DefaultValue :: * ;
import Assert       :: * ;
import Connectable  :: * ;

`include "Logger.bsv"
`include "trap.defines"

import pipe_ifcs    :: * ;
import dcache_types :: * ;
import csrbox       :: * ;
import csr_types    :: * ;
import ccore_types  :: * ;
import DReg         :: * ;

/*start*/

import bram         :: * ;

typedef 32 PC_WIDTH; // assuming 32-bit PC
typedef 10 TRACE_DEPTH; // 2^10 = 1024 entries

/*end*/

interface Ifc_stage5;
`ifdef debug
  interface Ifc_s5_debug debug;
`endif
`ifdef perfmonitors
  interface Ifc_s5_perfmonitors perf;
`endif
  interface Ifc_s5_rx rx;
  interface Ifc_s5_interrupts interrupts;
  interface Ifc_s5_common common;
  interface Ifc_s5_cache cache;
  interface Ifc_s5_csrs csrs;
endinterface:Ifc_stage5

/*start*/

UserInterface#(PC_WIDTH, PC_WIDTH, TAdd#(TRACE_DEPTH, 3)) trace_bram <- 
    mkbram(0, "trace_bram", "stage5");  // Set correct address base
Reg#(Bit#(TRACE_DEPTH)) trace_wr_ptr <- mkReg(0);

/*end*/

`ifdef stage5_noinline
/*doc:module: */
`ifdef core_clkgate
(*synthesize,gate_all_clocks*)
`else
(*synthesize*)
`endif
`endif
`ifdef simulate
(*preempts = "rl_writeback_memop, rl_no_op"*)
(*preempts = "rl_writeback_trap, rl_no_op"*)
(*preempts = "rl_writeback_system, rl_no_op"*)
(*preempts = "rl_writeback_baseout, rl_no_op"*)
`endif
module mkstage5#(parameter Bit#(`xlen) hartid) (Ifc_stage5);

  /*doc:submodules: The following instantiates all the RX virtual fifos*/
  RX#(SystemOut) rx_systemout <- mkRX;
  RX#(TrapOut)   rx_trapout <- mkRX;
  RX#(BaseOut)   rx_baseout <- mkRX;
  RX#(WBMemop)   rx_memio <- mkRX;
  RX#(CUid)      rx_fuid <- mkRX;
`ifdef rtldump
  RX#(CommitLogPacket) rx_commitlog <- mkRX;
`endif
 
  /*doc:submodules: The following instantiates the csr module generated by csrbox*/
  Ifc_csrbox csr <- mk_csrbox();

  /*doc:reg: This register holds the local epoch value of this stage*/
  Reg#(Bit#(1)) rg_epoch <- mkReg(0);

  /*doc:reg: This register when set is used to indicate that we need wait for the csrbox to respond*/
  Reg#(Bool) rg_csr_wait <- mkReg(False);

  /*doc:wire wire that carries the commit data that needs to be written to the integer register
   * file. IN cases of traps and instructions that need to be dropped, writing to this wire can be
   * used to release the lock on a register in the score-board*/
  Wire#(CommitData) wr_commit <- mkWire();

  /*doc:wire: This wire is used to indicate the rest of the pipeline that this stage has generated a
  * flush. In case of post-fenceI/sfence this signal also holds fields which are used to indicate
  * the I$ about a possible fenceI or sfence on the ITLB*/
  Wire#(WBFlush) wr_flush <- mkDWire(defaultValue);

  /*doc:wire: When set to True causes an increment in the minstret counter. Note in case of a csr
  * operation that writes a value to minstret. The new value of minstret at the end of the cycle
  * would be write-value + 1.*/
  Wire#(Bool) wr_increment_minstret <- mkDWire(False);

  /*doc:reg: This register when set indicates that an IO memory operation is in progress*/
  Reg#(Bool) rg_ioop_init <- mkReg(False);

  /*doc:wire: This wire holds the response of an IO memory operation */
  Wire#(Maybe#(DMem_core_response#(TMul#(`dwords,8),`desize))) wr_ioop_response <- mkDWire(tagged Invalid);

  /*doc:wire: this wire holds the epoch value of the IO memory store/atomic operation that is
   * waiting to be committed/dropped. Writing a value to this wire triggers an IO operation*/
  Wire#(Bit#(1)) wr_commit_ioop <- mkWire();

`ifdef dcache
  /*doc:wire: this wire holds the epoch value of the cached memory store/atomic operation that is
   * waiting to be committed/dropped*/
  Wire#(Tuple2#(Bit#(1), Bit#(TLog#(`dsbsize)))) wr_commit_cacheop <- mkWire();
`endif    
`ifdef debug
  /*doc:submodules: connection back to the csrs to stop counters*/
  mkConnection(csr.ma_stop_count, csr.mv_stop_count);
`endif
`ifdef rtldump
  /*doc:reg: When an instruction commits, this register holds the commit log packet in the next
   * cycle which can be consumed by the test-bench to write into a file*/
  Reg#(Maybe#(CommitLogPacket)) rg_commitlog <- mkDReg(tagged Invalid);
`endif
`ifdef perfmonitors
  /*doc:wire: wire to increment when exceptions detected*/
  Wire#(Bit#(1)) wr_count_exceptions <- mkDWire(0);
  /*doc:wire: wire to increment when interrupts detected*/
  Wire#(Bit#(1)) wr_count_interrupts <- mkDWire(0);
  /*doc:wire: wire to increment when csr-ops detected*/
  Wire#(Bit#(1)) wr_count_csrops <- mkDWire(0);
  /*doc:wire: wire to increment when micro-traps are detected*/
  Wire#(Bit#(1)) wr_count_microtrap <- mkDWire(0);
`endif

  let csr_response = csr.mv_core_resp;
  let epochs_match = rg_epoch == rx_fuid.u.first.epochs;

`ifdef simulate
  rule rl_no_op;
    `logLevel( stage5, 0, $format("[%2d]STAGE5: No Instr to commit", hartid))
  endrule: rl_no_op
`endif

  /*doc:rule: This rule handles all traps there were detected/raised in any of the previous stages
  * for any given instruction. The rule also checks if the micro-trap is generated and acts
  * accordingly. For a regular trap like load-access/load-page-fault, the load instruction would
  * have locked a register in the score-board and would thus require to be released inspite of
  * taking of the fault. To ensure this release, we update the wr_commit signal to make this release
  * on the destination register*/
  rule rl_writeback_trap(rx_fuid.u.first.insttype == TRAP );
    let trapout = rx_trapout.u.first;
    let fuid = rx_fuid.u.first;
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : PC:%h",hartid,fuid.pc))
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : Trap: ",hartid, fshow(trapout)))
    wr_commit <= CommitData{addr: fuid.rd, data: ?, unlock_only:True
                          `ifdef no_wawstalls , id: fuid.id `endif
                           `ifdef spfpu ,rdtype: fuid.rdtype `endif };

    if (epochs_match) begin
     /*start*/
     let pc = fuid.pc;
     trace_bram.write_request(tuple3(zeroExtend(trace_wr_ptr), pc, '1));
     trace_wr_ptr <= (trace_wr_ptr + 1) & ('h3FF);

     /*end*/

    `ifdef microtrap_support
      if (trapout.is_microtrap) begin
        if (trapout.cause == `Sfence_rerun || trapout.cause == `FenceI_rerun || 
            trapout.cause == `CSR_rerun 
					`ifdef hypervisor || trapout.cause == `Hfence_rerun `endif ) begin
          let _fencei = (trapout.cause == `FenceI_rerun);
          let _sfence = (trapout.cause == `Sfence_rerun);
  			  let _hfence = (trapout.cause == `Hfence_rerun);
          wr_flush <= WBFlush{flush: True, newpc : fuid.pc , fencei: _fencei 
              `ifdef supervisor , sfence: _sfence `endif 
              `ifdef hypervisor , hfence: _hfence `endif };
          `logLevel( stage5, 0, $format("[%2d]STAGE5 : Redirect PC:%h",hartid, fuid.pc))
        `ifdef perfmonitors
          wr_count_microtrap <= 1;
        `endif
        end
        else begin
          dynamicAssert(False, "Received unexpected Micro-Trap cause");
        end
      end
      else `endif begin
        let tvec <- csr.mav_upd_on_trap(trapout.cause, fuid.pc, trapout.mtval 
          `ifdef hypervisor , trapout.mtval2 `endif );
        wr_flush <= WBFlush{flush: True, newpc : tvec, fencei: False 
            `ifdef supervisor , sfence: False `endif 
            `ifdef hypervisor , hfence: False `endif };
      `ifdef perfmonitors
        Bit#(1) cause_type = truncateLSB(trapout.cause);
        if (cause_type == 1)
          wr_count_interrupts <= 1;
        else
          wr_count_exceptions <= 1;
      `endif
        `logLevel( stage5, 0, $format("[%2d]STAGE5 : Going to *TVEC:%h",hartid, tvec))
      end
        rx_trapout.u.deq;
        rx_fuid.u.deq;
        rg_epoch <= ~rg_epoch;
      `ifdef rtldump
        rx_commitlog.u.deq;
      `endif
    end
    else begin
      `logLevel( stage5, 0, $format("[%2d]STAGE5 : Dropping instruction",hartid))
      rx_trapout.u.deq;
      rx_fuid.u.deq;
    `ifdef rtldump
      rx_commitlog.u.deq;
    `endif
    end
  endrule:rl_writeback_trap

  /*doc:rule: This rule is used to commit system operations which could be xRET ops or CSR ops.
  * Committing a xRET ops causes a flush to be raised with a new pc coming from the csrbox. In case
  * of CSR ops, one might have to wait for multiple cycles for the execution to complete and then
  * commit the value.*/
  rule rl_writeback_system(rx_fuid.u.first.insttype == SYSTEM ) ;
    let systemout = rx_systemout.u.first;
    let fuid = rx_fuid.u.first;
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : PC:%h",hartid,fuid.pc))
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : ",hartid, fshow(systemout)))
    Bool exit = False;
    if (epochs_match) begin

      /*start*/
      let pc = fuid.pc;
      trace_bram.write_request(tuple3(zeroExtend(trace_wr_ptr), pc, '1));
      trace_wr_ptr <= (trace_wr_ptr + 1) & ('h3FF);

     /*end*/

      if (systemout.funct3 == 0 ) begin // URET, SRET, MRET
        let epc <- csr.mav_upd_on_ret(truncateLSB(systemout.csr_address));
        exit = True;
        wr_flush <= WBFlush{flush: True, newpc : epc, fencei: False
          `ifdef supervisor , sfence: False `endif 
          `ifdef hypervisor , hfence: False `endif };
        rg_epoch <= ~rg_epoch;
          `logLevel( stage5, 0, $format("[%2d]STAGE5 : Redirect PC:%h",hartid,epc))
      end
      else if (!rg_csr_wait) begin
        csr.ma_core_req(CSRReq{csr_address: systemout.csr_address, writedata: systemout.rs1_imm,
            funct3: truncate(systemout.funct3) `ifdef compressed , pc_1: fuid.pc[1] `endif });
      end
  
      if ((systemout.funct3 !=0 && csr_response.hit) || (systemout.funct3==0)) begin
        rg_csr_wait <= False;
        exit = True;
      end
      else begin
        rg_csr_wait <= True;
        `logLevel( stage5, 0, $format("[%2d]STAGE5 : Waiting for CSR-response",hartid))
      end
  
      if (exit) begin
        wr_increment_minstret <= True;
        wr_commit <= CommitData{addr: fuid.rd, data: zeroExtend(csr_response.data), unlock_only:False
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu ,rdtype: fuid.rdtype `endif };
        rx_systemout.u.deq;
        rx_fuid.u.deq;
      `ifdef perfmonitors
        if (systemout.funct3 != 0)
          wr_count_csrops <= 1;
      `endif
      `ifdef rtldump
        let clogpkt = rx_commitlog.u.first;
        CommitLogCSR _pkt = ?;
        if (clogpkt.inst_type matches tagged CSR .pcsr)
          _pkt = pcsr;
        if (systemout.funct3 == 0) begin
          _pkt.csr_address = 'h300;
          _pkt.wdata = csr.sbread.mv_csr_mstatus;
        end
        _pkt.rdata = csr_response.data;
        clogpkt.inst_type = tagged CSR _pkt;
        clogpkt.mode = csr.mv_prv;
			`ifdef hypervisor
				clogpkt.v = csr.mv_virtual;
			`endif
        rg_commitlog <= tagged Valid clogpkt;
        rx_commitlog.u.deq;
      `endif
      end
    end
    else begin
      `logLevel( stage5, 0, $format("[%2d]STAGE5 : Dropping instruction",hartid))
      wr_commit <= CommitData{addr: fuid.rd, data: ?, unlock_only:True
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu ,rdtype: fuid.rdtype `endif };
      rx_systemout.u.deq;
      rx_fuid.u.deq;
    `ifdef rtldump
      rx_commitlog.u.deq;
    `endif
    end
  endrule:rl_writeback_system

  /*doc:rule: This rule basically commits regular ops which update the register file. Note that even
  * Loads will land up here. So the commit log packet is not touched since it would be tagged
  * CommitLogMem for Loads which has to be passed on as is to the test-bench*/
  rule rl_writeback_baseout(rx_fuid.u.first.insttype == BASE);
    let fuid = rx_fuid.u.first;
    let baseout = rx_baseout.u.first;
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : PC:%h",hartid,rx_fuid.u.first.pc))
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : Base Op ",hartid, fshow(baseout)))
    if (epochs_match) begin
      wr_increment_minstret <= True;
      `ifdef spfpu csr.ma_set_fflags(baseout.fflags, fuid.rdtype); `endif
      wr_commit <= CommitData{addr: fuid.rd, data: zeroExtend(baseout.rdvalue), unlock_only:False
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu ,rdtype: fuid.rdtype `endif };
      /*start*/

      let pc = fuid.pc;
      trace_bram.write_request(tuple3(zeroExtend(trace_wr_ptr), pc, '1));
      trace_wr_ptr <= (trace_wr_ptr + 1) & ('h3FF);


      /*end*/
      rx_fuid.u.deq;
      rx_baseout.u.deq;
    `ifdef rtldump
      let clogpkt = rx_commitlog.u.first;
      rx_commitlog.u.deq;
      clogpkt.mode = csr.mv_prv;
			`ifdef hypervisor
				clogpkt.v = csr.mv_virtual;
			`endif
      rg_commitlog <= tagged Valid clogpkt;
    `endif
    end
    else begin
      `logLevel( stage5, 0, $format("[%2d]STAGE5 : Dropping instruction",hartid))
      wr_commit <= CommitData{addr: fuid.rd, data: ?, unlock_only:True
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu ,rdtype: fuid.rdtype `endif };
      rx_baseout.u.deq;
      rx_fuid.u.deq;
    `ifdef rtldump
      rx_commitlog.u.deq;
    `endif
    end
  endrule:rl_writeback_baseout

  /*doc:rule: This rule performs memory operations. In specific it completes a previously cached
  * store/atomic operation or initiates a new IO memory operation. This rule simply indicates the
  * Store buffer or the IO buffer held in the cache to initiate the respective operation. This
  * indication is basically a write to the wr_commit_cacheop/wr_commit_ioop wire with the current
  * epoch value.
  * In case a cached store/atomic op has to be dropped since the epochs don't match. The epoch value
  * sent will cause the respective entry in the caches to be dropped without any updates to cache/
  * memory*/
  rule rl_writeback_memop(rx_fuid.u.first.insttype == MEMORY );
    let memop = rx_memio.u.first;
    let fuid = rx_fuid.u.first;
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : PC:%h",hartid,fuid.pc))
  `ifdef rtldump
    let clogpkt = rx_commitlog.u.first;
    CommitLogMem _pkt = ?;
    if (clogpkt.inst_type matches tagged MEM. cmem) 
      _pkt = cmem;
  `endif

    if (epochs_match) begin

     /*start*/
     let pc = fuid.pc;
     trace_bram.write_request(tuple3(zeroExtend(trace_wr_ptr), pc, '1));
     trace_wr_ptr <= (trace_wr_ptr + 1) & ('h3FF);

     /*end*/

    `ifdef dcache
      if (!memop.io) begin // cacheable store/atomic op
        `logLevel( stage5, 0, $format("[%2d]STAGE5 : Cached Store Op ",hartid, fshow(memop)))
        wr_commit_cacheop <= tuple2(rg_epoch, memop.sb_id);
        wr_increment_minstret <= True;
        rx_fuid.u.deq;
        rx_memio.u.deq;
      `ifdef atomic
        let cache_resp = memop.atomic_rd_data;
        if (memop.memaccess == Atomic) 
          wr_commit <= CommitData{addr: fuid.rd, data: zeroExtend(cache_resp), unlock_only:False
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu ,rdtype: fuid.rdtype `endif };
      `else
        Bit#(`elen) cache_resp = 0;
      `endif
      `ifdef rtldump
        rx_commitlog.u.deq;
        _pkt.commit_data = cache_resp;
        clogpkt.inst_type = tagged MEM _pkt;
        clogpkt.mode = csr.mv_prv;
			`ifdef hypervisor
				clogpkt.v = csr.mv_virtual;
			`endif
        rg_commitlog <= tagged Valid clogpkt;
      `endif
      end
      else 
    `endif
      begin 
        `logLevel( stage5, 0, $format("[%2d]STAGE5 : Non-Cached Memory Op ",hartid, fshow(memop)))
        if (!rg_ioop_init) begin
          rg_ioop_init <= True;
          wr_commit_ioop <= rg_epoch;
        end
        else if (wr_ioop_response matches tagged Valid .ioresp) begin
          rg_ioop_init <= False;
          if (ioresp.trap) begin
            let tvec <- csr.mav_upd_on_trap(ioresp.cause, fuid.pc, ioresp.word 
            `ifdef hypervisor , ? `endif 
            );
            wr_flush <= WBFlush{flush: True, newpc : tvec, fencei: False 
                `ifdef supervisor , sfence: False `endif 
                `ifdef hypervisor , hfence: False `endif };
            `logLevel( stage5, 0, $format("[%2d]STAGE5 : Redirect PC:%h",hartid, tvec))
            rg_epoch <= ~rg_epoch;
            rx_fuid.u.deq;
            rx_memio.u.deq;
            wr_commit <= CommitData{addr: fuid.rd, data: ?, unlock_only: True
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu ,rdtype: fuid.rdtype `endif };
          `ifdef rtldump
            rx_commitlog.u.deq;
          `endif
          end
          else begin
            wr_increment_minstret <= True;
            let commit_data = ioresp.word;
            `ifdef dpfpu if (memop.nanboxing) commit_data[63:32] = '1; `endif
            wr_commit <= CommitData{addr: fuid.rd, data: zeroExtend(commit_data), unlock_only:False
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu ,rdtype: fuid.rdtype `endif };
            rx_fuid.u.deq;
            rx_memio.u.deq;
          `ifdef rtldump
            rx_commitlog.u.deq;
            _pkt.commit_data = (fuid.rd ==0 `ifdef spfpu && fuid.rdtype == IRF `endif )?0:commit_data;
            clogpkt.inst_type = tagged MEM _pkt;
            clogpkt.mode = csr.mv_prv;
					`ifdef hypervisor
						clogpkt.v = csr.mv_virtual;
					`endif
            rg_commitlog <= tagged Valid clogpkt;
          `endif
          end
        end
        else begin
          `logLevel( stage5, 0, $format("[%2d]STAGE5: Waiting for IO response",hartid))
        end
      end
    end
    else begin
      `logLevel( stage5, 0, $format("[%2d]STAGE5 : Dropping instruction",hartid))
      wr_commit <= CommitData{addr: fuid.rd, data: ?, unlock_only:True
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu ,rdtype: fuid.rdtype `endif };
      rx_memio.u.deq;
      rx_fuid.u.deq;
    `ifdef rtldump
      rx_commitlog.u.deq;
    `endif
    `ifdef dcache
      if(!memop.io)
        wr_commit_cacheop <= tuple2(rg_epoch, ?);
      else
    `endif
        wr_commit_ioop <= rg_epoch;
    end
  endrule:rl_writeback_memop

  /*doc:rule: This rule is fired when wr_increment_minstret is set and thus cases the minstret
  * register to increment*/
  rule rl_incr_minstret(wr_increment_minstret);
    csr.ma_incr_minstret(1);
  endrule:rl_incr_minstret

  interface rx = interface Ifc_s5_rx
    interface rx_systemout_from_stage4  = rx_systemout.e;
    interface rx_trapout_from_stage4  = rx_trapout.e;
    interface rx_baseout_from_stage4 = rx_baseout.e;
    interface rx_memio_from_stage4 = rx_memio.e;
    interface rx_fuid_from_stage4 = rx_fuid.e;
  `ifdef rtldump
    interface rx_commitlog = rx_commitlog.e;
  `endif
  endinterface;
  
  interface interrupts = interface Ifc_s5_interrupts
    method ma_clint_msip = csr.ma_set_mip_msip;
    method ma_clint_mtip = csr.ma_set_mip_mtip;
    // if time register is not needed, then mtime value is not required
    // time register is used in user mode
    `ifdef user
    method ma_clint_mtime = csr.ma_set_time;
    `endif
    method ma_plic_meip = csr.ma_set_mip_meip;
  `ifdef hypervisor
  	method ma_plic_vseip = csr.ma_set_vseip;
  `endif
  `ifdef supervisor 
    method ma_plic_seip = csr.ma_set_mip_seip;
  `endif
  `ifdef usertraps
    method ma_plic_ueip = csr.ma_set_mip_ueip;
  `endif
  endinterface;
`ifdef debug 
  interface debug = interface Ifc_s5_debug
    method mv_csr_dcsr = csr.sbread.mv_csr_dcsr;
    method ma_debug_interrupt= csr.ma_set_mip_debug_interrupt;
    method mv_debug_mode= csr.mv_debug_mode;
    method mv_core_debugenable = csr.sbread.mv_csr_customcontrol[4];
    method mv_stop_timer = csr.mv_stop_timer;
    method mv_stop_count = csr.mv_stop_count;
  endinterface;
`endif

`ifdef perfmonitors
  interface perf = interface Ifc_s5_perfmonitors
    method ma_events = csr.ma_events;
   	method mv_count_exceptions = wr_count_exceptions;
   	method mv_count_interrupts = wr_count_interrupts;
   	method mv_count_csrops = wr_count_csrops;
   	method mv_count_microtraps = wr_count_microtrap;
  endinterface;
`endif
  
  interface common = interface Ifc_s5_common
    method mv_commit_rd = wr_commit;
    method mv_flush = wr_flush;
  `ifdef rtldump
    method mv_commit_log = rg_commitlog;
  `endif
  endinterface;
  
  interface cache = interface Ifc_s5_cache
    method mv_initiate_store = wr_commit_cacheop;
    method Bit#(1) mv_initiate_ioop = wr_commit_ioop;
    method Action ma_io_response(Maybe#(DMem_core_response#(TMul#(`dwords,8),`desize)) r);
      wr_ioop_response <= r;
    endmethod:ma_io_response
  endinterface;
  interface csrs = interface Ifc_s5_csrs;
    method mv_csr_misa_c = csr.sbread.mv_csr_misa[2];
    method mv_cacheenable = truncate(csr.sbread.mv_csr_customcontrol);
    method mv_curr_priv = pack(csr.mv_prv);
    method mv_csr_mstatus = csr.sbread.mv_csr_mstatus;
  `ifdef hypervisor
		`ifdef RV32
			method mv_csr_mstatush = csr.sbread.mv_csr_mstatush;
 		`endif
		method mv_csr_hstatus = csr.sbread.mv_csr_hstatus;
		method mv_csr_vsstatus = csr.sbread.mv_csr_vsstatus;				
		method mv_csr_vsatp = csr.sbread.mv_csr_vsatp;
		method mv_csr_hgatp = csr.sbread.mv_csr_hgatp;
		method mv_vs_bit = csr.mv_virtual;
  `endif
    method mv_csrs_to_decode = CSRtoDecode {prv: csr.mv_prv,
        csr_mip: truncate(csr.sbread.mv_csr_mip), 
        csr_mie: truncate(csr.sbread.mv_csr_mie), 
        csr_mstatus: truncate(csr.sbread.mv_csr_mstatus),
        csr_sstatus: `ifdef hypervisor (csr.mv_virtual == 1)? csr.sbread.mv_csr_vsstatus: `endif csr.sbread.mv_csr_mstatus,
        csr_misa: truncate(csr.sbread.mv_csr_misa)
      `ifdef spfpu
        ,frm: truncate(csr.sbread.mv_csr_frm)
      `endif
      `ifdef debug
        ,csr_dcsr: truncate(csr.sbread.mv_csr_dcsr)
      `endif
      `ifdef non_m_traps 
        ,csr_mideleg: truncate(csr.sbread.mv_csr_mideleg)
    `endif 
    `ifdef hypervisor
    , csr_hideleg: truncate(csr.sbread.mv_csr_hideleg)
    , csr_hstatus: truncate(csr.sbread.mv_csr_hstatus)   
    , csr_vs_bit: truncate(csr.mv_virtual)
      `endif };
    method mv_resume_wfi = unpack( |((csr.sbread.mv_csr_mip)& (csr.sbread.mv_csr_mie) ));
	`ifdef supervisor
		method mv_csr_satp = csr.sbread.mv_csr_satp;
	`endif
  `ifdef pmp
    method mv_pmp_cfg = csr.mv_pmpcfg;
    method mv_pmp_addr = csr.mv_pmpaddr;
  `endif
  `ifdef rtldump
    interface sbread = csr.sbread;
  `endif
  endinterface;
endmodule: mkstage5

endpackage: stage5

Sdram.bsv:

/* 
Copyright (c) 2018, IIT Madras All rights reserved.

Redistribution and use in source and binary forms, with or without modification, are permitted
provided that the following conditions are met:

* Redistributions of source code must retain the above copyright notice, this list of conditions
  and the following disclaimer.  
* Redistributions in binary form must reproduce the above copyright notice, this list of 
  conditions and the following disclaimer in the documentation and/or other materials provided 
 with the distribution.  
* Neither the name of IIT Madras nor the names of its contributors may be used to endorse or 
  promote products derived from this software without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS
OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, 
DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER
IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT 
OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--------------------------------------------------------------------------------------------------

Copyright (c) 2018, IIT Madras All rights reserved.

Redistribution and use in source and binary forms, with or without modification, are permitted
provided that the following conditions are met:

* Redistributions of source code must retain the above copyright notice, this list of conditions
  and the following disclaimer.  
* Redistributions in binary form must reproduce the above copyright notice, this list of 
  conditions and the following disclaimer in the documentation and/or other materials provided 
 with the distribution.  
* Neither the name of IIT Madras  nor the names of its contributors may be used to endorse or 
  promote products derived from this software without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS
OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER
IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT 
OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--------------------------------------------------------------------------------------------------
*/


package sdram;
`include "sdram.defines"
import Semi_FIFOF        :: *;
import AXI4_Types   :: *;
import AXI4_Fabric  :: *;
import bsvmksdrc_top :: *;
import BUtils            ::*;
import Connectable ::*;
import ConfigReg ::*;
import DReg::*;
import FIFOF::*;
import Clocks::*;
import device_common::*;

/*start*/
import bram :: *;
typedef 32 PC_WIDTH; // assuming 32-bit PC
typedef 10 TRACE_DEPTH; // 2^10 = 1024 entries

parameter Integer TRACE_BRAM_BASE = 32'h9000_0000;
Ifc_bram_axi4#(PC_WIDTH, 0, PC_WIDTH, 0, TAdd#(TRACE_DEPTH, 3)) ifc_trace_bram_axi4 <- mkbram_axi4(TRACE_BRAM_BASE, "trace_bram") clocked_by clk0 reset_by rst0;
/*end*/

export Ifc_sdram_out      (..);
export Ifc_sdram_axi4     (..); // interface export
export mksdram_axi4;        // module export  

/*start*/
export Ifc_trace_bram_axi4(..);
interface Ifc_trace_bram_axi4;
    interface AXI4_Slave_IFC#(PC_WIDTH, 0, PC_WIDTH, 0) slave_trace_bram;
endinterface

interface trace_bram_axi4 = ifc_trace_bram_axi4.slave;
/*end*/
  

interface Ifc_sdram_out#(numeric type io_width);
	(*always_enabled,always_ready*)
    method Action ipad_sdr_din(Bit#(io_width) pad_sdr_din);
    method Bit#(9) sdram_sdio_ctrl();
    method Bit#(io_width) osdr_dout();
    method Bit#(8) osdr_den_n();
    method Bool osdr_cke();
    method Bool osdr_cs_n();
    method Bool osdr_ras_n ();
    method Bool osdr_cas_n ();
    method Bool osdr_we_n ();
    method Bit#(8) osdr_dqm ();
    method Bit#(2) osdr_ba ();
    method Bit#(13) osdr_addr ();
    interface Clock sdram_clk;    
endinterface

interface Ifc_sdram_axi4#(numeric type addr_width, 
                           numeric type data_width, 
                           numeric type user_width,
                           numeric type io_width,
                           numeric type rfrsh_timer_width,
                           numeric type rfrsh_row_width);                       
      interface AXI4_Slave_IFC#(addr_width, data_width, user_width) slave_mem;
      interface AXI4_Slave_IFC#(addr_width, data_width, user_width) slave_cfg;
      interface Ifc_sdram_out#(io_width) io;
endinterface

typedef enum{
    IDLE,
    WRITE_START,
    WAIT_DELAY,
    WRITE_FIRST,
    WRITE_DATA0,
    WRITE_DATA1
} Write_state deriving(Bits, Eq, FShow);

typedef enum{
    IDLE,
    START_READ,
    READ_DATA,
    READ_FLUSH
} Read_state deriving(Bits, Eq,FShow);

typedef enum {
    IDLE,
    START_SPLIT,
    SEND_VALUE
} Write_split_states deriving(Bits, Eq, FShow);


function (Bit#(9)) fn_wr_len(Bit#(8) length, Bit#(3) awsize, Bit#(3) lwr_addr);
     Bit#(3) w_packet = 0;
     Bit#(9) s_length = 0;
 case(awsize)
        
     'd0 : begin
         w_packet = lwr_addr >> awsize;
         s_length = ((zeroExtend(length) + zeroExtend(w_packet)) >> 3) + 1;
     end
     'd1: begin
         w_packet = lwr_addr >> awsize;
         s_length = ((zeroExtend(length) + zeroExtend(w_packet)) >> 2) + 1;
 //`ifdef verbose $display($time(),"\t SSSS w_packet %b s_lenght %h length %h", w_packet, s_length, length); `endif
     end
     'd2 : begin
        //w_packet = lwr_addr >> awsize;
        // s_length = ((s_length + w_packets) >> 1) + 1;
        s_length = zeroExtend(length >> 1) + 1;
     end
     'd3 : begin
         s_length = zeroExtend(length) + 1;
     end
 endcase

 return s_length;
endfunction


function Bit#(26) fn_wr_address(Bit#(addr_width) address);
    Bit#(29) sdr_addr = address[31:3];
    return sdr_addr[25:0];
endfunction




//(*synthesize*)
    
module mksdram_axi4#(Clock clk0, Reset rst0) (Ifc_sdram_axi4#(addr_width, 
                                                      data_width, 
                                                      user_width,
                                                      io_width,
                                                      rfrsh_timer_width,
                                                      rfrsh_row_width))
                                                      provisos(
                                                         Add#(e__, 1, data_width),
                                                         Add#(g__, 2, data_width),
                                                         Add#(h__, 3, data_width),
                                                         Add#(i__, 4, data_width),
                                                         Add#(f__, 13, data_width),
                                                         Add#(a__, 8, data_width),
                                                         Add#(b__, 9, data_width),
                                                         Add#(c__, 12, data_width),
                                                         Add#(d__, 8, addr_width),
                                                         Add#(j__, data_width, 64),
                                                        Mul#(strb, 8, data_width),
                                                        Div#(data_width, 8, strb),
                                                Add#(k__, 8, TDiv#(data_width, 8)),
                                                Add#(l__, rfrsh_row_width, data_width),
                                                Add#(m__, rfrsh_timer_width, data_width),
                                                Add#(n__, 3, rfrsh_row_width),
                                                Add#(o__, 12, rfrsh_timer_width),
//                                                SizedLiteral#(Bit#(rfrsh_timer_width), 12),
//                                                SizedLiteral#(Bit#(rfrsh_row_width), 3),
                                                Add#(p__, data_width, io_width),
                                                Add#(q__, io_width, data_width)
                                                      );
    
function Bit#(data_width) fn_wr_split_data(Bit#(data_width) data, Bit#(strb) wstrb);
    Bit#(data_width) data0 = 0;
    Bit#(8) temp_data0 = 0;
    for(Integer i=0; i<valueOf(strb); i=i+1) begin
        if(wstrb[i]==1)
            temp_data0 = data[8*(i)+7:8*(i)];
            data0[8*(i)+7:8*(i)] = temp_data0; 
    end
//    if(wstrb[0] == 1)
//        data0[7:0] = data[7:0];
//    else
//        data0[7:0] = 0;
//
//    if(wstrb[1] == 1)
//        data0[15:8] = data[15:8];
//    else
//        data0[15:8] = 0;
//
//    if(wstrb[2] == 1)
//        data0[23:16] = data[23:16];
//    else
//        data0[23:16] = 0;
//
//    if(wstrb[3] == 1)
//        data0[31:24] = data[31:24];
//    else
//        data0[31:24] = 0;
//
//    if(wstrb[4] == 1)
//        data0[39:32] = data[39:32];
//    else
//        data0[39:32] = 0;
//
//    if(wstrb[5] == 1)
//        data0[47:40] = data[47:40];
//    else
//        data0[47:40] = 0;
//
//    if(wstrb[6] == 1)
//        data0[55:48] = data[55:48];
//    else
//        data0[55:48] = 0;
//
//    if(wstrb[7] == 1)
//        data0[63:56] = data[63:56];
//    else
//        data0[63:56] = 0;
//
    return data0;
endfunction

function Bit#(data_width) fn_rd_data(Bit#(3) bsize,Bit#(6) lwr_addr,Bit#(data_width) data);
    //Integer b_strb = valueOf(TLog#(strb));
    Bit#(64) max_width=0;
    Bit#(64) in_data = zeroExtend(data);
    if(bsize=='b000) begin
        Bit#(8) out_data = in_data[((8) * (lwr_addr+1)) - 1 : (8 * lwr_addr)];
        max_width = duplicate(out_data);
    end
    if(bsize=='b001) begin
        Bit#(16) out_data = in_data[((16) * (lwr_addr+1)) - 1 : (16 * lwr_addr)];
        max_width = duplicate(out_data);
    end
    if(bsize=='b010) begin
        Bit#(32) out_data = in_data[((32) * (lwr_addr+1)) - 1 : (32 * lwr_addr)];
        max_width = duplicate(out_data);
    end
    if(valueOf(data_width)==64) begin
        if(bsize=='b011) begin
            Bit#(64) out_data = in_data; 
            max_width = out_data;
        end
    end
    return truncate(max_width);
//    case(bsize)
//        'b000: begin
//            case(lwr_addr)
//                'b000: begin
//                    max_width = duplicate(data[7:0]);
//                end
//                'b001: begin
//                    max_width = duplicate(data[15:8]);
//                end
//                'b010: begin
//                    max_width = duplicate(data[23:16]);
//                end
//                'b011: begin
//                    max_width = duplicate(data[31:24]);
//                end
//                'b100: begin
//                    max_width = duplicate(data[39:32]);
//                end
//                'b101: begin
//                    max_width = duplicate(data[47:40]);
//                end
//                'b110: begin
//                    max_width = duplicate(data[55:48]);
//                end
//                'b111: begin
//                    max_width = duplicate(data[63:56]);
//                end
//            endcase
//        end
//
//        'b001: begin
//    return duplicate(data[lwr_addr[b_strb*16] : lwr_addr[(bstrb-1)*16]])
//            case(lwr_addr) 
//                'b000: begin
//                    max_width = duplicate(data[15:0]);
//                end
//                'b010: begin
//                    max_width = duplicate(data[31:16]);
//                end
//                'b100: begin
//                    max_width = duplicate(data[47:32]);
//                end
//                'b110: begin
//                    max_width = duplicate(data[63:48]);
//                end
//            endcase
//        end
//
//        'b010: begin
//            case(lwr_addr)
//                'b000: begin
//                    max_width = duplicate(data[31:0]);
//                end
//                'b100: begin
//                    max_width = duplicate(data[63:32]);
//                end
//            endcase
//        end
//        'b011: begin
//            if(valueOf(data_width)==64)
//                max_width = data;
//        end
//    endcase
//    return truncate(max_width);
endfunction

//Reset rst0 <- mkAsyncResetFromCR (0, clk0);

Reg#(Bit#(9))        rg_delay_count <- mkRegA(0,clocked_by clk0, reset_by rst0);
Reg#(Bit#(9))        rg_rd_actual_len <- mkRegA(0,clocked_by clk0, reset_by rst0);
Reg#(bit)            rg_app_req <- mkDRegA(0,clocked_by clk0, reset_by rst0);
Reg#(bit)            rg_app_req_wrap <- mkConfigRegA(0,clocked_by clk0, reset_by rst0);
Reg#(Bit#(26))       rg_app_req_addr <- mkConfigRegA(0,clocked_by clk0, reset_by rst0);
Reg#(Bit#(4))        rg_cfg_sdr_tras_d <- mkConfigRegA(4'h4,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(4))        rg_cfg_sdr_trp_d <- mkConfigRegA(4'h2,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(4))        rg_cfg_sdr_trcd_d <- mkConfigRegA(4'h2,clocked_by clk0, reset_by rst0); 
Reg#(bit)            rg_cfg_sdr_en <- mkConfigRegA(1'h0,clocked_by clk0, reset_by rst0);
Reg#(Bit#(2))        rg_cfg_req_depth <- mkConfigRegA(2'h3,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(13))       rg_cfg_sdr_mode_reg <- mkConfigRegA(13'h032,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(3))        rg_cfg_sdr_cas <- mkConfigRegA(3'h3,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(4))        rg_cfg_sdr_trcar_d <- mkConfigRegA(4'h7,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(4))        rg_cfg_sdr_twr_d <- mkConfigRegA(4'h1,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(2))        rg_cfg_sdr_width <- mkConfigRegA(2'b0,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(2))        rg_cfg_colbits <- mkConfigRegA(2'b01,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(9))        rg_cfg_sdio_ctrl <- mkConfigRegA(9'b000100011,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(8))        rg_cfg_sdr_clk_delay <- mkConfigRegA(8'b00001000,clocked_by clk0, reset_by rst0);

Reg#(Bit#(rfrsh_timer_width ))  rg_cfg_sdr_rfsh <- mkConfigRegA('h100,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(rfrsh_row_width)) rg_cfg_sdr_rfmax <- mkConfigRegA('h6,clocked_by clk0, reset_by rst0); 
Reg#(Bit#(9))                   rg_app_req_len <- mkConfigRegA(0,clocked_by clk0, reset_by rst0);
Reg#(Bit#(4))                   rg_lwraddr <- mkConfigRegA(0,clocked_by clk0, reset_by rst0);
Reg#(Bit#(3))                   rg_arsize <- mkConfigRegA(0,clocked_by clk0, reset_by rst0);
Reg#(bit)                       rg_app_req_wr_n <- mkConfigRegA(0,clocked_by clk0, reset_by rst0);
Reg#(Bit#(TDiv#(data_width,8)))                   rg_app_wr_en_n <- mkDWire('hFF,clocked_by clk0, reset_by rst0);
Reg#(Bit#(data_width))                  rg_app_wr_data <- mkDWire(0,clocked_by clk0, reset_by rst0);
Wire#(Bool)                     wr_sdr_init_done <- mkDWire(False,clocked_by clk0, reset_by rst0);
Wire#(Bool)                     wr_app_req_ack <- mkDWire(False,clocked_by clk0, reset_by rst0);
Wire#(Bool)                     wr_app_wr_next_req <- mkDWire(False,clocked_by clk0, reset_by rst0);
Wire#(Bool)                     wr_app_rd_valid <- mkDWire(False,clocked_by clk0, reset_by rst0);
Wire#(Bool)                     wr_app_last_rd <- mkDWire(False,clocked_by clk0, reset_by rst0);
Wire#(Bool)                     wr_app_last_wr <- mkDWire(False,clocked_by clk0, reset_by rst0);
Wire#(Bit#(data_width))                 wr_app_rd_data <- mkWire(clocked_by clk0, reset_by rst0);


Reg#(Bit#(4))     rg_rid          <- mkRegA(0, clocked_by clk0, reset_by rst0);
Reg#(bit)         rg_rd_not_active_flag <- mkSyncRegToCC(0,clk0, rst0);
Reg#(Bit#(4))     rg_ctrl_rid     <- mkRegA(0);
Reg#(Bit#(4))     rg_wid          <- mkRegA(0);

Reg#(Write_split_states) rg_wr_split_states <- mkRegA(IDLE); 
Reg#(Bit#(3))            rg_awsize          <- mkRegA(0);
Reg#(Bit#(9))            rg_ac_count        <- mkRegA(0);
Reg#(Bit#(6))            rg_single_burst    <- mkRegA(0);
Reg#(Bit#(data_width))           rg_wr_ac_data      <- mkRegA(0);
Reg#(Bit#(TDiv#(data_width,8)))            rg_wr_ac_wstrb     <- mkRegA(0);
Reg#(Bit#(4))            rg_wr_lwr_addr     <- mkRegA(0); 
Reg#(Bit#(9))            rg_local_actual_wr_length <- mkRegA(0);
Reg#(Bit#(9))            rg_actual_wr_length <- mkSyncRegFromCC(0,clk0);
Reg#(Bit#(addr_width))           rg_wr_address       <- mkSyncRegFromCC(0,clk0);

Reg#(Bit#(3))            rg_awsize_sclk       <- mkSyncRegFromCC(0,clk0);

Reg#(Bit#(9))            rg_burst_counter        <- mkRegA(0);

Bool burst_eq = (rg_burst_counter == rg_local_actual_wr_length);

Reg#(Bit#(3))          rg_packets          <- mkRegA(0);
Reg#(Bit#(3))          rg_packet_counter   <- mkRegA(0);


Reg#(Write_state) rg_write_states <- mkRegA(IDLE,clocked_by clk0, reset_by rst0);
Reg#(Read_state) rg_read_states <- mkRegA(IDLE,clocked_by clk0, reset_by rst0);

FIFOF#(AXI4_Wr_Addr#(addr_width, user_width)) ff_wr_addr        <- mkSizedFIFOF(13);
FIFOF#(AXI4_Wr_Data#(data_width))        ff_wr_data        <- mkSizedFIFOF(13);
SyncFIFOIfc#(Bit#(data_width))           ff_ac_wr_data     <- mkSyncFIFOFromCC(13,clk0);
SyncFIFOIfc#(Bit#(TDiv#(data_width,8)))                    ff_ac_wr_wstrb    <- mkSyncFIFOFromCC(13,clk0);

SyncFIFOIfc#(Bool) ff_sync_write_response<-mkSyncFIFOToCC(1,clk0,rst0);

   //FIFOF#(AXI4_Rd_Addr#(addr_width,user_width)) ff_rd_addr <- mkSizedFIFOF(3);
FIFOF#(Bit#(data_width)) ff_rd_data <- mkSizedFIFOF(86,clocked_by clk0, reset_by rst0);
SyncFIFOIfc#(AXI4_Rd_Addr#(addr_width, user_width)) ff_rd_addr <- mkSyncFIFOFromCC(30,clk0);
SyncFIFOIfc#(AXI4_Rd_Data#(data_width, user_width)) ff_sync_read_response <-mkSyncFIFOToCC(13,clk0,rst0);

SyncFIFOIfc#(Tuple2#(Bit#(addr_width),Bit#(data_width))) ff_sync_ctrl_write<- mkSyncFIFOFromCC(1,clk0);
SyncFIFOIfc#(Bit#(addr_width)) ff_sync_ctrl_read<- mkSyncFIFOFromCC(1,clk0);
SyncFIFOIfc#(Bit#(data_width)) ff_sync_ctrl_read_response<- mkSyncFIFOToCC(1,clk0,rst0);

// Polling Registers
Reg#(Bit#(2)) rg_poll_cnt <- mkRegA(0,clocked_by clk0, reset_by rst0);
Reg#(Bool)    rg_polling_status <- mkSyncRegToCC(False,clk0,rst0);
Reg#(Bool)    rg_polling_status_clk0 <- mkRegA(False,clocked_by clk0, reset_by rst0);
Reg#(Bool)    rg_rd_trnc_flg <- mkRegA(False);
Reg#(Bool)    rg_wr_trnc_flg <- mkRegA(False);
Reg#(bit)     rg_odd_len     <- mkRegA(0);   
// hardcoding the parameter value to resolve provisos
AXI4_Slave_Xactor_IFC #(addr_width, data_width, user_width)  s_xactor_sdram     <- mkAXI4_Slave_Xactor;
AXI4_Slave_Xactor_IFC #(addr_width, data_width, user_width)  s_xactor_cntrl_reg <- mkAXI4_Slave_Xactor;
Ifc_sdram#(io_width, rfrsh_timer_width, rfrsh_row_width) sdr_cntrl <- mksdrc_top(clocked_by clk0, reset_by rst0);

function Action fn_wr_cntrl_reg(Bit#(data_width) data, Bit#(addr_width) address);
   
   action
   Bit#(8) addr = truncate(address);
   case(truncate(addr)) 

       `ACTPRE_DELAY    : rg_cfg_sdr_tras_d <= data[3:0];

       `PREACT_DELAY    : rg_cfg_sdr_trp_d <= data[3:0];
       
       `ACT_RW_DELAY    : rg_cfg_sdr_trcd_d <= data[3:0];
      
       `EN_SDRAM        : rg_cfg_sdr_en <= data[0];
      
       `MAX_REQ         : rg_cfg_req_depth <= data[1:0];
      
       `MODE_REG        : rg_cfg_sdr_mode_reg <= data[12:0];
      
       `CAS_LATNCY      : rg_cfg_sdr_cas <= data[2:0];
      
       `AUTO_REFRESH    : rg_cfg_sdr_trcar_d <= data[3:0];
      
       `RECRY_DELAY     : rg_cfg_sdr_twr_d <= data[3:0];
     // 
       `RFRSH_TIMER     : rg_cfg_sdr_rfsh <= extend(data[11:0]);

       `RFRSH_ROW_CNT   : rg_cfg_sdr_rfmax <= extend(data[2:0]);

       `SDR_WIDTH       : rg_cfg_sdr_width <= data [1:0];

       `SDR_COLBITS     : rg_cfg_colbits <= data [1:0];
       
       `SDR_SDIO_CTRL   : rg_cfg_sdio_ctrl <= data [8:0];

       `SDR_CLK_DELAY   : rg_cfg_sdr_clk_delay <= data [7:0];

       default          : noAction;
  endcase
  endaction 
endfunction

function Bit#(data_width) fn_rd_cntrl_reg(Bit#(addr_width) address);
//    provisos(
//             Add#(a__, 1, data_width),
//             Add#(b__, 2, data_width),
//             Add#(c__, 8, data_width),
//             Add#(d__, 9, data_width),
//             Add#(e__, 12, data_width),
//             Add#(f__, 13, data_width),
//             Add#(g__, 8, addr_width)
//            );
  Bit#(8) addr = truncate(address);
  case(addr)

       `ACTPRE_DELAY    :  return extend(rg_cfg_sdr_tras_d);

       `PREACT_DELAY    :  return extend(rg_cfg_sdr_trp_d);
       
       `ACT_RW_DELAY    :  return extend(rg_cfg_sdr_trcd_d);
      
       `EN_SDRAM        :  return extend(rg_cfg_sdr_en);
      
       `MAX_REQ         :  return extend(rg_cfg_req_depth);
      
       `MODE_REG        :  return extend(rg_cfg_sdr_mode_reg);
      
       `CAS_LATNCY      :  return extend(rg_cfg_sdr_cas);
      
       `AUTO_REFRESH    :  return extend(rg_cfg_sdr_trcar_d);
      
       `RECRY_DELAY     : return extend(rg_cfg_sdr_twr_d);
      
       `RFRSH_TIMER     : return extend(rg_cfg_sdr_rfsh);

       `RFRSH_ROW_CNT   : return extend(rg_cfg_sdr_rfmax);

       `SDR_INIT_DONE   : return extend(pack(wr_sdr_init_done));

       `SDR_WIDTH       : return extend(rg_cfg_sdr_width);

       `SDR_COLBITS     : return extend(rg_cfg_colbits);

       `SDR_SDIO_CTRL   : return extend(rg_cfg_sdio_ctrl);

       `SDR_CLK_DELAY   : return extend(rg_cfg_sdr_clk_delay);

    endcase 
endfunction
          
//(*preempts="(rl_pop_read_request, rl_send_rd_data, rl_send_read_data, rl_flush_redundant_data), rl_write_transaction_write_start"*)

rule rl_for_writing_ctrl_reg(ff_sync_ctrl_write.notFull);
    let aw <- pop_o(s_xactor_cntrl_reg.o_wr_addr);
    let w  <- pop_o(s_xactor_cntrl_reg.o_wr_data);
    `ifdef verbose $display($time,"\tSDRAM: control_reg written addr %x data %x", aw.awaddr, w.wdata); `endif
	  ff_sync_ctrl_write.enq(tuple2(aw.awaddr,w.wdata));
    let w_resp = AXI4_Wr_Resp {bresp: AXI4_OKAY, buser: 0, bid: aw.awid}; 
    s_xactor_cntrl_reg.i_wr_resp.enq(w_resp);
endrule

rule rl_perform_write_to_ctrl(ff_sync_ctrl_write.notEmpty);
	let {awaddr,wdata}=ff_sync_ctrl_write.first;
  `ifdef verbose $display("\tSDRAM: "); `endif
	ff_sync_ctrl_write.deq;
`ifdef verbose $display($time,"\tSDRAM: Actually writing data: %h to addr: %h", wdata, awaddr); `endif
    fn_wr_cntrl_reg(wdata , truncate(awaddr));    
endrule

rule rl_for_read_cntrl_reg;
    let ar <- pop_o(s_xactor_cntrl_reg.o_rd_addr);
	  ff_sync_ctrl_read.enq(ar.araddr);
	  rg_ctrl_rid<=ar.arid;
 endrule

 rule rl_send_ctrl_read_response(ff_sync_ctrl_read.notEmpty);
	 ff_sync_ctrl_read_response.enq(fn_rd_cntrl_reg(truncate(ff_sync_ctrl_read.first)));
	 ff_sync_ctrl_read.deq;
endrule

rule sync_ctr_response(ff_sync_ctrl_read_response.notEmpty);
	ff_sync_ctrl_read_response.deq;
    let r = AXI4_Rd_Data {rresp: AXI4_OKAY, rdata:ff_sync_ctrl_read_response.first ,
    rlast: True, ruser: 0, rid: rg_ctrl_rid};
    s_xactor_cntrl_reg.i_rd_data.enq(r);
endrule

rule rl_direct_connection_insdram;
    sdr_cntrl.iapp_req(rg_app_req);
    sdr_cntrl.iapp_req_wrap(rg_app_req_wrap);
    sdr_cntrl.iapp_req_addr(rg_app_req_addr);
    sdr_cntrl.iapp_req_len(rg_app_req_len);
    sdr_cntrl.iapp_req_wr_n(rg_app_req_wr_n);
    sdr_cntrl.iapp_wr_data(extend(rg_app_wr_data));
    sdr_cntrl.iapp_wr_en_n(truncate(rg_app_wr_en_n));
endrule

rule rl_direct_connection_outsdram;
    wr_sdr_init_done <= sdr_cntrl.osdr_init_done ;
    wr_app_req_ack <= sdr_cntrl.oapp_req_ack ();
    wr_app_wr_next_req <= sdr_cntrl.oapp_wr_next_req ();
    wr_app_rd_valid <= sdr_cntrl.oapp_rd_valid ();
    wr_app_last_rd <= sdr_cntrl.oapp_last_rd ();
    wr_app_last_wr <= sdr_cntrl.oapp_last_wr ();
    wr_app_rd_data <= extend(sdr_cntrl.oapp_rd_data);
endrule

rule rl_direct_connection_config_reg;
    sdr_cntrl.icfg_sdr_tras_d(rg_cfg_sdr_tras_d);
    sdr_cntrl.icfg_sdr_trp_d(rg_cfg_sdr_trp_d);
    sdr_cntrl.icfg_sdr_trcd_d(rg_cfg_sdr_trcd_d);
    sdr_cntrl.icfg_sdr_en(rg_cfg_sdr_en);
    sdr_cntrl.icfg_req_depth(rg_cfg_req_depth);
    sdr_cntrl.icfg_sdr_mode_reg(rg_cfg_sdr_mode_reg);
    sdr_cntrl.icfg_sdr_cas(rg_cfg_sdr_cas);
    sdr_cntrl.icfg_sdr_trcar_d(rg_cfg_sdr_trcar_d);
    sdr_cntrl.icfg_sdr_twr_d(rg_cfg_sdr_twr_d);
    sdr_cntrl.icfg_sdr_rfsh(rg_cfg_sdr_rfsh);
    sdr_cntrl.icfg_sdr_rfmax(rg_cfg_sdr_rfmax);
    sdr_cntrl.icfg_sdr_width(rg_cfg_sdr_width);
    sdr_cntrl.icfg_colbits(rg_cfg_colbits);
endrule

rule rl_intial_polling(rg_polling_status_clk0 == False && wr_sdr_init_done == True);
    `ifdef verbose	$display($time,"\tSDRAM: POLLING MODE: %d",rg_poll_cnt); `endif 
    case (rg_poll_cnt)
        0: begin
            rg_app_req <= 1;
            rg_app_req_addr <= 0;
            rg_app_req_len <= 1;
            rg_app_req_wr_n <= 0;
            rg_app_wr_en_n <= 'hFF;
            rg_app_wr_data <= 0;
            rg_poll_cnt <= rg_poll_cnt + 1;
        end
        1: begin
            rg_app_req <= 1;
            rg_app_req_addr <= 0;
            rg_app_req_len <= 1;
            rg_app_req_wr_n <= 0;
            rg_app_wr_en_n <= 'hFF;
            rg_app_wr_data <= 0;
            rg_poll_cnt <= rg_poll_cnt + 1;
        end
        2: begin
            rg_app_req <= 0;
            rg_app_req_addr <= 0;
            rg_app_wr_en_n <= 'hFF;
            rg_app_wr_data <= 0;
            if(wr_app_wr_next_req == True)
                rg_poll_cnt <= rg_poll_cnt + 1;
        end
        3: begin
            rg_polling_status <= True;
				 rg_polling_status_clk0<=True;
        end
    endcase
endrule

/******************* WRITE TRANSACTION ****************/

rule rl_parallel_data_enq(rg_polling_status == True && rg_rd_trnc_flg == False);
    let aw <- pop_o(s_xactor_sdram.o_wr_addr);
    let w  <- pop_o(s_xactor_sdram.o_wr_data);
    ff_wr_addr.enq(aw);
    ff_wr_data.enq(w);      
    rg_wr_trnc_flg <= True;
    `ifdef verbose $display($time,"\tSDRAM: WRITE_FIRST Parallel enq %h addr: %h",w.wdata,aw.awaddr); `endif
endrule

rule rl_write_split_state(rg_wr_split_states == IDLE);
    let aw = ff_wr_addr.first();
    if(aw.awsize != 3) begin
        rg_actual_wr_length <= fn_wr_len(aw.awlen, aw.awsize, aw.awaddr[2:0]);

        rg_local_actual_wr_length <= extend(aw.awlen);
    end
    else begin
        rg_actual_wr_length <= extend(aw.awlen) + 1;
        rg_local_actual_wr_length <= extend(aw.awlen);
    end
    rg_wid <= aw.awid;
    rg_awsize <= aw.awsize;
    rg_awsize_sclk <= aw.awsize;
    rg_wr_address <= aw.awaddr;
    rg_wr_lwr_addr <= extend(aw.awaddr[2:0]);
    rg_wr_split_states <= START_SPLIT;
    rg_packets <=  (aw.awsize==0)?7:(aw.awsize==1)?3:(aw.awsize == 2)? 1 : (aw.awsize == 3) ? 0 : 0; //(64 >> (aw.awsize+4));  //1 << ~aw.awsize[1:0];
    rg_packet_counter <= (aw.awaddr[2:0]) >> aw.awsize;
    `ifdef verbose $display($time,"Initial Values -- Starting IDLE to START_SPLIT"); `endif
    //$display("Initial Values: rg_packets: %h rg_packet_counter: %h ",(64>>(aw.awsize+4)),aw.awaddr[2:0]>>aw.awsize);
    rg_burst_counter <= 0;
endrule


rule rl_write_data_splitting0(rg_wr_split_states == START_SPLIT && rg_awsize != 3);
   rg_wr_ac_data <= rg_wr_ac_data | fn_wr_split_data(ff_wr_data.first.wdata,ff_wr_data.first.wstrb);
   rg_wr_ac_wstrb <= rg_wr_ac_wstrb | ff_wr_data.first.wstrb;
   rg_burst_counter <= rg_burst_counter + 1;
   //`ifdef verbose $display($time,"burst_eq: %h rg_packets: %h rg_packet_counter: %d rg_burst_counter: %d rg_local_actual_wr_length %d rg_wr_ac_data %h rg_wr_ac_wstrb %b",burst_eq,rg_packets,rg_packet_counter
   //,rg_burst_counter,rg_local_actual_wr_length, fn_wr_split_data(ff_wr_data.first.wdata,ff_wr_data.first.wstrb),
   //ff_wr_data.first.wstrb); `endif
       if(burst_eq || rg_packets == rg_packet_counter) begin
           rg_wr_split_states <= SEND_VALUE;
       end
       else begin
          rg_packet_counter <= rg_packet_counter + 1;
       end
        ff_wr_data.deq();
        ff_wr_addr.deq();
endrule

rule rl_write_data_splitting1(rg_wr_split_states == SEND_VALUE && rg_awsize != 3);
    `ifdef verbose $display($stime,"Splitting1 Enqueued data rg_wr_ac_data %h rg_wr_ac_wstrb %b", rg_wr_ac_data, rg_wr_ac_wstrb); `endif
    ff_ac_wr_data.enq(rg_wr_ac_data);
    ff_ac_wr_wstrb.enq(rg_wr_ac_wstrb);
    rg_wr_ac_data <= 0;            
    rg_wr_ac_wstrb <= 0;
    rg_wr_lwr_addr <= 0;
    rg_packet_counter <= 0;
    `ifdef verbose $display($time,"Sending Value to the SDRAM"); `endif
    rg_wr_split_states <= START_SPLIT;
endrule

rule rl_write_data_spliting3(rg_wr_split_states == START_SPLIT && rg_awsize == 3);
    ff_ac_wr_data.enq(ff_wr_data.first.wdata);
    ff_ac_wr_wstrb.enq(ff_wr_data.first.wstrb);
    ff_wr_data.deq();
    ff_wr_addr.deq();
endrule

rule rl_start_write_transaction(rg_write_states == IDLE && wr_sdr_init_done == True);        
    if(ff_ac_wr_data.notEmpty()) begin
        if(rg_awsize_sclk == 0)
            rg_write_states <= WAIT_DELAY;
        else
        rg_write_states <= WRITE_START;
        `ifdef verbose $display($time,"\tSDRAM: Going to write start state"); `endif
    end
endrule

rule rl_wait_delay(rg_write_states == WAIT_DELAY);
    if(rg_delay_count == 14) begin
        rg_write_states <= WRITE_START;
        rg_delay_count <= 0;
    end
    else
    rg_delay_count <= rg_delay_count + 1;
endrule

rule rl_write_transaction_write_start(rg_write_states == WRITE_START && wr_sdr_init_done == True && rg_read_states == IDLE);
    `ifdef verbose $display($time,"\tSDRAM: WRITE_START state Controller Length %d",rg_actual_wr_length); `endif
    rg_app_req <= 1;
    rg_app_req_addr <= fn_wr_address(rg_wr_address);
    rg_app_req_len <= extend(rg_actual_wr_length);
    rg_app_req_wr_n <= 0;
    rg_app_wr_data <= 0;
    rg_app_wr_en_n <= 'hFF;
    rg_write_states <= WRITE_FIRST;
    rg_delay_count <= extend(rg_actual_wr_length) - 1;
endrule

rule rl_write_transaction_write_first(rg_write_states == WRITE_FIRST && wr_app_wr_next_req == False);
    `ifdef verbose $display($time,"\tSDRAM: WRITE_FIRST state next is false data %x",ff_ac_wr_data.first); `endif
    rg_app_req <= 0;
    rg_app_wr_en_n <= ~(ff_ac_wr_wstrb.first());
    rg_app_wr_data <= ff_ac_wr_data.first();               
endrule

rule rl_write_transaction_write_data(rg_write_states == WRITE_FIRST && wr_app_wr_next_req == True);
`ifdef verbose $display($time,"\tSDRAM: WRITE_DATA state next is true sending data %x %b",ff_ac_wr_data.first,
wr_app_wr_next_req); `endif
    rg_app_req <= 0;
    rg_app_wr_data <= ff_ac_wr_data.first();
    rg_app_wr_en_n <= ~(ff_ac_wr_wstrb.first());
    ff_ac_wr_data.deq;
    ff_ac_wr_wstrb.deq;
    rg_delay_count <= rg_delay_count - 1;
    if(rg_delay_count == 0) begin
       rg_write_states <= IDLE;
			ff_sync_write_response.enq(True);
    end
endrule

rule synchronize_write_response(ff_sync_write_response.notEmpty);
	ff_sync_write_response.deq;
	let w_resp = AXI4_Wr_Resp {bresp: AXI4_OKAY, buser: 0, bid: rg_wid}; //TODO user value is null
  s_xactor_sdram.i_wr_resp.enq(w_resp);
   rg_wr_split_states <= IDLE;
   rg_ac_count <= 0;
   rg_wr_trnc_flg <= False;
  `ifdef verbose   $display($time,"\tSDRAM: WRITE complete state true"); `endif
endrule
    
   /****************** Read Transaction ********************/
	//	`ifdef verbose
	//	  rule display_read_states;
	//		$display($time,"\tSDRAM: Read State: ",fshow(rg_read_states));
	//	  endrule
	//	`endif
rule rl_paralel_read_req_enq(rg_polling_status == True && rg_wr_trnc_flg == False);
    let ar <- pop_o(s_xactor_sdram.o_rd_addr);
     ff_rd_addr.enq(ar);
     rg_rd_trnc_flg <= True;
    `ifdef verbose	$display($time,"\tSDRAM: Got Read request from AXI for AddresS: %h",ar.araddr); `endif
endrule

rule rl_read_idle_state(rg_read_states == IDLE);
    if(ff_rd_addr.notEmpty() == True) begin
        rg_read_states <= START_READ;
        rg_rd_not_active_flag <= 0;
        `ifdef verbose  $display($time,"\tSDRAM: READ IDLE state"); `endif
    end

endrule

rule rl_pop_read_request(wr_sdr_init_done == True && rg_read_states == START_READ && (rg_write_states == IDLE || 
rg_write_states == WRITE_START));
let ar = ff_rd_addr.first;
`ifdef verbose $display($time,"\tSDRAM: STAR_READ state ar.arlen %d ar.arsize %d ar.araddr %h ar.arburst %b", ar.
arlen,ar.arsize, ar.araddr, ar.arburst); `endif

rg_app_req <= 1;
if(ar.arburst == 2)
    rg_app_req_wrap <= 1;
else
    rg_app_req_wrap <= 0;
rg_lwraddr <= extend(ar.araddr[2:0]);
rg_arsize <= ar.arsize;
rg_app_req_addr <= fn_wr_address(ar.araddr);
rg_app_req_len <= fn_wr_len(ar.arlen, ar.arsize, ar.araddr[2:0]);
rg_rd_actual_len <= extend(ar.arlen);
rg_app_req_wr_n <= 1;
rg_delay_count <= 0;
rg_read_states <= READ_DATA;
rg_rid <= ar.arid;
`ifdef verbose $display($time,"\t SSSSS SDRAM START_READ length "); `endif
endrule

rule rl_send_rd_data(wr_app_rd_valid == True);
    `ifdef verbose $display($time,"\tSDRAM: READ DATA1 state %x",wr_app_rd_data); `endif
    ff_rd_data.enq(wr_app_rd_data);
endrule

rule rl_send_read_data(rg_read_states==READ_DATA);
`ifdef verbose $display($time,"\tSDRAM: Response from BFM. RequestLenght: %d CurrentCount: %d",rg_rd_actual_len,
rg_delay_count); `endif
rg_app_req_wrap <= 0;
if(rg_lwraddr < 8) begin
      let r = AXI4_Rd_Data {rresp: AXI4_OKAY, rdata: fn_rd_data(rg_arsize, extend(rg_lwraddr), ff_rd_data.first), rlast: 
      (rg_rd_actual_len == rg_delay_count), ruser: 0, rid: rg_rid};
  		  ff_sync_read_response.enq(r);
  		  ff_rd_addr.deq;
  		  if(rg_arsize!=3)
          rg_lwraddr <= rg_lwraddr + (1 << rg_arsize);
  			else
  				ff_rd_data.deq;
  		//`ifdef verbose $display($time,"\tSDRAM: SENDING READ DATA : %h, rg_lwraddr %b rg_arsize %d", 
         // fn_rd_data(rg_arsize, rg_lwraddr, ff_rd_data.first),rg_lwraddr, rg_arsize); `endif
  			`ifdef verbose $display($time,"\tSDRAM: Removing Request for Addr : %h",ff_rd_addr.first.araddr); `endif
   if(rg_delay_count == rg_rd_actual_len) begin
    `ifdef verbose  $display($time,"\tSDRAM: SENT ALL READ DATA state rg_delay_count %d rg_rd_actual_len %d", 
    rg_delay_count, rg_rd_actual_len); `endif
      rg_read_states <= READ_FLUSH;
      rg_rd_not_active_flag <= 1;
      rg_delay_count <= 0;
   end
   else 
     rg_delay_count <= rg_delay_count + 1;
 end
 else if(rg_lwraddr > 7) begin
        `ifdef verbose $display($time,"\tSDRAM: Dequeuing ff READ"); `endif
        rg_lwraddr <= 0;
        ff_rd_data.deq;
 end
endrule

rule rl_flush_redundant_data(rg_read_states == READ_FLUSH);
    ff_rd_data.clear();
    rg_read_states <= IDLE;
endrule

rule send_synchronized_read_response(ff_sync_read_response.notEmpty);
  let r=ff_sync_read_response.first;
  `ifdef verbose	$display($time,"\tSDRAM: Sending Read response: %h rlast: %b",r.rdata,r.rlast); `endif
  ff_sync_read_response.deq;
  if(rg_rd_not_active_flag == 1)
  rg_rd_trnc_flg <= False;
  s_xactor_sdram.i_rd_data.enq(r);
endrule


interface Ifc_sdram_out io;

    method Action ipad_sdr_din(Bit#(io_width) pad_sdr_din);
        sdr_cntrl.ipad_sdr_din(pad_sdr_din);
    endmethod
    method Bit#(9) sdram_sdio_ctrl();
        return rg_cfg_sdio_ctrl;
    endmethod
    method Bit#(io_width) osdr_dout();
        return sdr_cntrl.osdr_dout();
    endmethod
    method Bit#(8) osdr_den_n();
        return sdr_cntrl.osdr_den_n();
    endmethod
    method Bool osdr_cke();
        return sdr_cntrl.osdr_cke();
    endmethod

    method Bool osdr_cs_n();
        return sdr_cntrl.osdr_cs_n();
    endmethod

    method Bool osdr_ras_n ();
        return sdr_cntrl.osdr_ras_n;
    endmethod

    method Bool osdr_cas_n ();
        return sdr_cntrl.osdr_cas_n;
    endmethod

    method Bool osdr_we_n ();
        return sdr_cntrl.osdr_we_n;
    endmethod

    method Bit#(8) osdr_dqm ();
        return sdr_cntrl.osdr_dqm;
    endmethod

    method Bit#(2) osdr_ba ();
        return sdr_cntrl.osdr_ba;
    endmethod

    method Bit#(13) osdr_addr ();
        return sdr_cntrl.osdr_addr;
    endmethod
    
    interface sdram_clk = clk0;
endinterface
interface slave_mem= s_xactor_sdram.axi_side;
interface slave_cfg = s_xactor_cntrl_reg.axi_side;

endmodule
endpackage
Ccore.bsv:

// See LICENSE.iitm for license details
/*

Author : IIT Madras
Details:

--------------------------------------------------------------------------------------------------
*/
package ccore;

//=================== Interface and module for a ccore - master on the AXI4 fabric ============= //
// project related imports
import Semi_FIFOF:: *;
import AXI4_Types:: *;
import AXI4_Fabric:: *;
//import riscv:: * ;
import riscv :: *;
import ccore_types:: * ;
import FIFOF::*;
import dcache_types :: *;
import icache_types :: * ;
import Assert ::*;
import imem::*;
import dmem::*;
import pipe_ifcs :: * ;
/*start*/
import sdram :: *;
import bram  :: *;
typedef 32 PC_WIDTH; // assuming 32-bit PC
typedef 10 TRACE_DEPTH; // 2^10 = 1024 entries

/*end*/
`ifdef hypervisor
  import ptwalk_hypervisor :: * ;
`elsif supervisor
  import ptwalk_merged::*;
`endif
`include "ccore_params.defines"
`include "Logger.bsv"


`define Mem_master_num 0

// package imports
import Connectable 				:: *;
import GetPut:: *;
import BUtils::*;
import csrbox :: * ;

`ifdef debug
import debug_types  :: * ;
import csr_types    :: * ;
`endif

`ifdef supervisor
typedef enum {None, IWalk, DWalk} PTWState deriving(Bits, Eq, FShow);
`endif

interface Ifc_ccore_axi4;
	interface AXI4_Master_IFC#(`paddr, `axi4_id_width, `buswidth, USERSPACE) master_d;
	interface AXI4_Master_IFC#(`paddr, `axi4_id_width, `buswidth, USERSPACE) master_i;
    interface Put#(Bit#(1)) sb_clint_msip;

	/*doc:method: This method should receive the machine timer interrupt from the CLINT module*/
  interface Put#(Bit#(1)) sb_clint_mtip;

	/*doc:method: This method should receive the machine timer value from the CLINT module. This will
	* be used for the pseduo op rdtime instruction in the user mode*/
  interface Put#(Bit#(64)) sb_clint_mtime;

  /*doc:method: This method should receive the machine external interrupt from the PLIC module*/
	method Action sb_plic_meip(Bit#(1) ex_i);

`ifdef supervisor
  /*doc:method: When supervisor is enabled, this method will receive the supervisor external
   * interrupt from the PLIC. Note this is a different context from the machine external interrupt*/
	method Action sb_plic_seip(Bit#(1) ex_i);
`endif
`ifdef usertraps
  /*doc:method: When user traps (N-extesion) is enabled, this method will receive the user external
   * interrupt from the PLIC. Note this is a different context from the machine,supervisor 
   * external interrupt*/
	method Action sb_plic_ueip(Bit#(1) ex_i);
`endif
`ifdef rtldump
  /*doc:sbifc: This interface is available only for simulation when intruction trace dump has been 
  enabled. This method is used to read the value of the csrs in the next cycle after csr-ops are
  done. This allows the TB to dump the correct value that is written to the csr.*/
  interface Sbread sbread;
  /*doc:method: this method carries the trace dump information of the instruction that was recently
   * committed*/
  method Maybe#(CommitLogPacket) commitlog;
`endif
`ifdef debug
  /*doc:method: This method is used to capture the interrupt from the debugger in case of resume or
   * halt indication*/
  method Action ma_debug_interrupt(Bit#(1) _int);
  /*doc:method: This method indicates if the core has been reset successfully*/
  method Bit#(1) mv_core_is_reset;

  /*doc:method: This method indicates to the debugger is the core is available for debugging*/
  method Bit#(1) mv_core_debugenable;

`ifndef core_clkgate
  (*always_enabled*)
`endif
  /*doc:method: This action method indicates the core that a debugger is connected and available for
   * carrying our debug operations*/
  method Action ma_debugger_available (Bit#(1) avail);
  /*doc:method: This method holds the bits from the dcsr register which indicate that the timer in
   * CLINT should stop incrementing when in debug mode*/
  method Bit#(1) mv_stop_timer;
  /*doc:method: This method holds the bits from the dcsr register which indicate that the
   * mhpmcounters in the csrs should stop incrementing when in debug mode*/
  method Bit#(1) mv_stop_count;
`endif
endinterface : Ifc_ccore_axi4

`ifdef core_clkgate
  (*synthesize,gate_all_clocks*)
`else
  (*synthesize*)
`endif
`ifdef supervisor
  (*preempts="rl_dtlb_req_to_ptwalk, rl_itlb_req_to_ptwalk"*)
  (*preempts="core_req_mkConnectionGetPut, ptwalk_req_mkConnectionGetPut"*)
`endif

`ifdef itim
  (*conflict_free="handle_itim_write_resp, handle_nc_write_resp"*)
`endif
(*mutually_exclusive ="rl_handle_io_read_response, rl_handle_io_write_resp"*)
module mkccore_axi4#(Bit#(`vaddr) resetpc, parameter Bit#(`xlen) hartid `ifdef testmode ,Bool test_mode `endif )(Ifc_ccore_axi4);
  String core = "";
  /*doc:mod: instatiate the riscv pipeline */
  
  /*start*/
  parameter Integer SDRAM_BASE = 32'h80000000;
  parameter Integer SDRAM_SIZE = 32'h10000000;
  parameter Integer TRACE_BRAM_BASE = 32'h90000000;
  parameter Integer TRACE_BRAM_SIZE = 32'h00001000;

  /*end*/

  Ifc_riscv riscv <- mkriscv(resetpc, hartid `ifdef testmode ,test_mode `endif );

  /*start*/
  Ifc_sdram_axi4 sdram <- mksdram_axi4(...);
  Ifc_trace_bram_axi4 trace_bram <- mkbram_axi4(TRACE_BRAM_BASE, "trace_bram");

  function Bit#(1) addr_decode (Bit#(32) addr);
        if ((addr >= SDRAM_BASE) && (addr < SDRAM_BASE+SDRAM_SIZE)) return 0;
        else if ((addr >= TRACE_BRAM_BASE) && (addr < TRACE_BRAM_BASE+TRACE_BRAM_SIZE)) return 1;
        else return 0; // default/fault/error
    endfunction
  /*end*/

  `ifdef supervisor
    Reg#(PTWState) rg_ptw_state <- mkReg(None);
  `endif
    `ifdef hypervisor
    Ifc_ptwalk ptwalk <- mkptwalk;
  `elsif supervisor
    Ifc_ptwalk#(`asidwidth) ptwalk <- mkptwalk;
  `endif

	AXI4_Master_Xactor_IFC #(`paddr, `axi4_id_width , `buswidth, USERSPACE) fetch_xactor <- mkAXI4_Master_Xactor;
	AXI4_Master_Xactor_IFC #(`paddr, `axi4_id_width ,`buswidth, USERSPACE) memory_xactor <- mkAXI4_Master_Xactor;
        /*start*/
        AXI4_Fabric_IFC #(NUM_MASTERS, 2, 32, ID_WIDTH, 32, USER_WIDTH) fabric <- mkAXI4_Fabric(addr_decode);

 fabric.v_to_slaves = vector(sdram.slave_mem, trace_bram.slave_trace_bram);
 fabric.v_from_masters = vector(fetch_xactor.axi_side, memory_xactor.axi_side);

       /*end*/

`ifdef pmp
  /*doc:var: When pmp is enabled we capture the curernt pmp configurations and addresses that will
  * be required by the TLBs*/
  let lv_pmp_cfg = riscv.csrs.mv_pmp_cfg;
  let lv_pmp_adr = riscv.csrs.mv_pmp_addr;
`endif

  /*doc:mod: instantiate the instruction memory subsystem*/
	Ifc_imem imem <- mkimem(truncate(hartid) `ifdef pmp ,lv_pmp_cfg, lv_pmp_adr `endif  `ifdef testmode ,test_mode `endif );

  /*doc:mod: instantiate the data memory subsystem*/
	Ifc_dmem dmem <- mkdmem(truncate(hartid) `ifdef pmp ,lv_pmp_cfg, lv_pmp_adr `endif  `ifdef testmode ,test_mode `endif );

`ifdef dcache
  /*doc:reg: This register is used to keep track of the beats/bursts occurring during the write
  * operation of a data line to memory. A new line-write or an io-write operation can be initiated
  * only when rg_burst_count == 0, else the requests are stalled. */
  Reg#(Bit#(8)) rg_burst_count <- mkReg(0);

  /*doc:reg: While performing burst writes during line eviction, this register indicates the amount
   * the line should be shifted to send the next beat of data on the bus*/
  Reg#(Bit#(TLog#(TMul#(TMul#(`dwords, 8), `dblocks)))) rg_shift_amount <- mkReg(`buswidth);
`endif
  /*doc: capture the current privilege mode under which the current transaction is being carried
  * out. TODO: This should ideally come form the caches themselves. Capturing here can have issues.
  * For example during an eviction, if the prv changes in the write-back stage then stores of the same
  * line may occur in different privilege modes*/
  let curr_priv = riscv.csrs.mv_curr_priv;

	/*doc:connect: Connect the instruction request from the core to the instruction memory subsystem*/
	mkConnection(imem.put_core_req , riscv.s0_icache.to_icache);

  /*doc:connect: Connect the instruction memory subsystem's response to the pipeline's stage-1 which
   * will accept it and process*/
	mkConnection(imem.get_core_resp, riscv.s1_icache.inst_response); // imem integration

  /*doc:connect: Send the signal from the data memory subsystem indicating that it is available to
   * receive new instructions from the stage3. If unavailable, stage3 should stall on a possible
   * memory operation.*/
	mkConnection(dmem.mv_dmem_available, riscv.s3_cache.ma_cache_is_available);

  /*doc:connect: Connect the load/store request happening in the stage3 of the pipeline to the
   * request port of the data memory subsystem*/
  let core_req <- mkConnection(dmem.receive_core_req, riscv.s3_cache.mv_memory_request);

  /*doc:connect: Connect the data memory subsystem's response to stage4 of the pipeline*/
	let core_resp <- mkConnection(dmem.send_core_cache_resp, riscv.s4_cache.memory_response); // dmem integration

  /*doc:rule: This rule sends out requests from the I-cache to the fabric. This rule will only fire
  * when there has been a line-miss in the instructino cache or the request is an io operation. This
  * rule also will not fire if the fetch-xactor fifo is full - which can happen due to contention in
  * the fabric*/
  rule rl_handle_imem_line_request;
		let request <- imem.get_read_mem_req.get;
		AXI4_Rd_Addr#(`paddr,`axi4_id_width, 0) imem_request = AXI4_Rd_Addr {araddr : truncate(request.address),
      aruser: ?, arlen : request.burst_len, arsize : request.burst_size, arburst : 'b10,
      arid : zeroExtend(pack(request.io)), arprot:{1'b1, 1'b0, curr_priv[1]} }; // arburst : 00 - FIXED 01 - INCR 10 - WRAP
	  fetch_xactor.i_rd_addr.enq(imem_request);
		`logLevel( core, 1, $format("[%2d]CORE : IMEM Line Requesting ",hartid, fshow(imem_request)))
  endrule:rl_handle_imem_line_request

  /*doc:rule: This rule captures the response from the fetch transactor of the fabric and routes
   * the response back to the instruction memory subsystem. This rule will fire only when the
   * fetch-xactor has a response available. The instruction memory is implicitly assumed to be always
   * available to pick the responses owing to its blocking nature*/
	rule rl_handle_imem_line_resp;
	  let fab_resp <- pop_o (fetch_xactor.o_rd_data);
		Bool bus_error = !(fab_resp.rresp == AXI4_OKAY);
    imem.put_read_mem_resp.put(ICache_mem_readresp{data   : truncate(fab_resp.rdata),
                                               last   : fab_resp.rlast,
                                               err    : bus_error,
                                               io     : (fab_resp.rid==1)});
		`logLevel( core, 1, $format("[%2d]CORE : IMEM Line Response ",hartid, fshow(fab_resp)))
	endrule:rl_handle_imem_line_resp

`ifdef icache
  /*doc:rule: This rule is used connect the cache enable signal for the instruction memory
   * subsystem*/
  rule rl_imem_enable;
	  imem.ma_cache_enable(unpack(riscv.csrs.mv_cacheenable[0]));
  endrule: rl_imem_enable
`endif

`ifdef dtim
  /*doc:rule: */
  rule rl_connect_dtim_memorymap_csrs;
    dmem.ma_dtim_memory_map(truncate(riscv.mv_csr_dtim_base), truncate(riscv.mv_csr_dtim_bound));
  endrule
`endif
`ifdef itim
  /*doc:rule: */
  rule rl_connect_itim_memorymap_csrs;
    imem.ma_itim_memory_map(truncate(riscv.mv_csr_itim_base), truncate(riscv.mv_csr_itim_bound));
  endrule
`endif

	/*doc:rule: This rule will initiate an IO read or write as indicated by the WB stage of the
	* pipeline. If a burst write is on-going then this rule is stalled. Since AXI4 support narrow
  * transfers (transfers whose size is lesser than the size of the bus), for write operations 
  * we make sure to duplicate
  * the data accordingly so that respective bytes of the lane contain the correct data. This is easier
  * than to shift the data.*/
  rule rl_initiate_io `ifdef dcache (rg_burst_count == 0) `endif ;
	  // receive the request from the data memory subsystem
	  let req <- dmem.send_mem_io_req.get;
    `logLevel( core, 0, $format("CORE: Received io op: ",fshow(req)))

    // resize the data and duplicate the bytes based on the size of the transaction 
   if(req.size[1:0]== 0)
      req.data = duplicate(req.data[7 : 0]);
    else if(req.size[1:0] == 1)
      req.data = duplicate(req.data[15 : 0]);
    else if(req.size[1:0] == 2)
      req.data = duplicate(req.data[31 : 0]);
     else 
       req.data = duplicate(req.data[63 : 0]);

    // build the write-strobe based on the size of the request.
    Bit#(TDiv#(`buswidth, 8)) write_strobe = req.size[1:0] == 0?'b1 :
                                        req.size[1:0] == 1?'b11 :
                                        req.size[1:0] == 2?'hf : 
                                        req.size[1:0] == 3?'hff :   '1;
    Bit#(TAdd#(1, TDiv#(`buswidth, 32))) byte_offset = truncate(req.address);
    write_strobe = write_strobe<<byte_offset;

    // if read operation send transaction on the i_rd_addr channel
	  if (!req.read_write) begin
		  AXI4_Rd_Addr#(`paddr,`axi4_id_width, 0) dmem_request = AXI4_Rd_Addr {araddr : truncate(req.address), aruser: ?,
        arlen : 0, arsize : zeroExtend(req.size[1:0]), arburst : 'b00, // arburst : 00 - FIXED 01 - INCR 10 - WRAP
        arid : 1 ,arprot:{1'b0, 1'b0, curr_priv[1]} }; 
      memory_xactor.i_rd_addr.enq(dmem_request);
	  end
	  // if write operation send transaction on the i_wr_addr and i_wr_data channels
	  else begin
	    AXI4_Wr_Addr#(`paddr,`axi4_id_width, 0) aw = AXI4_Wr_Addr {awaddr : truncate(req.address), awuser : 0,
        awlen : 0, awsize : zeroExtend(req.size[1 : 0]), awburst : 'b0,
        awid : 1, awprot:{1'b0, 1'b0, curr_priv[1]} }; // arburst : 00 - FIXED 01 - INCR 10 - WRAP

	let w  = AXI4_Wr_Data {wdata : truncate(req.data), wstrb : write_strobe,
                             wlast : True, 
                             wid : 1};
	    memory_xactor.i_wr_addr.enq(aw);
	    memory_xactor.i_wr_data.enq(w);
	  end
	endrule:rl_initiate_io

   /*doc:rule: This rule will receive the response generated for a previous data memory subsystem IO
  * read transaction. Because of the in-order nature of the core and that all IO transactions in the
  * WB stage can only be initiated when the previous one is over, we do not need to handle the
  * scenario where the responses can be out of order.*/
  rule rl_handle_io_read_response(memory_xactor.o_rd_data.first.rid == 1);
    let response <- pop_o(memory_xactor.o_rd_data);
  	let bus_error = !(response.rresp == AXI4_OKAY);
    dmem.receive_mem_io_resp.put(DCache_io_response{data:truncate(response.rdata), 
                                              error:bus_error});
    `logLevel( core, 1, $format("[%2d]CORE : IO Read Response ",hartid, fshow(response)))
  endrule:rl_handle_io_read_response


  /*doc:rule: This rule will receive the response generated for a previous data memory subsystem IO
  * write transaction. Because of the in-order nature of the core and that all IO transactions in the
  * WB stage can only be initiated when the previous one is over, we do not need to handle the
  * scenario where the responses can be out of order.*/
  rule rl_handle_io_write_resp (memory_xactor.o_wr_resp.first.bid == 1);
    let response <- pop_o(memory_xactor.o_wr_resp);
  	let bus_error = !(response.bresp == AXI4_OKAY);
    dmem.receive_mem_io_resp.put(DCache_io_response{data: ?, 
                                              error:bus_error});
    `logLevel( core, 1, $format("[%2d]CORE : IO Write Response ",hartid, fshow(response)))
  endrule:rl_handle_io_write_resp

`ifdef dcache

  /*doc:reg: This register when Valid, indicaets that there is pending read line operation which got
   * delayed because of a contentious write happening on the same line address*/
  Reg#(Maybe#(AXI4_Rd_Addr#(`paddr,`axi4_id_width, 0))) rg_read_line_req <- mkReg(tagged Invalid);

  /*doc:reg: This register when Valid, indicates the address to which a line a request is in
   * progress. This is used to delay a read operation on the same line initiated by the cache*/
  Reg#(Maybe#(Bit#(`paddr))) wr_write_req <- mkReg(tagged Invalid);
  
  /*doc:rule: This rule is used connect the cache enable signal for the data memory
   * subsystem*/
  rule rl_map_dmem_enable;
	  dmem.ma_cache_enable(unpack(riscv.csrs.mv_cacheenable[1]));
  endrule:rl_map_dmem_enable

  /*doc:connect: This connects the store commit routine from the WB stage of the pipeline to the
   * commit store method of the data memory subsystem*/
  mkConnection(dmem.ma_commit_store, riscv.s5_cache.mv_initiate_store);

  /*doc:connect: This connects the IO commit routine from the WB stage of the pipeline to the
   * commit io method of the data memory subsystem*/
  mkConnection(dmem.ma_commit_io, riscv.s5_cache.mv_initiate_ioop);

  /*doc:connect: This connects the io response from the data memory subsystem to the WB stage of the
   * pipeline */
  mkConnection(dmem.send_core_io_resp, riscv.s5_cache.ma_io_response);

  /*doc:rule: Currently it is possible that the data cache can generate a write - request followed by a
  read - request, but the fabric (due to contention) latches the read first to the slave followed
  by the write - req. This could lead to wrong behavior. To avoid this it is necessary to ensure
  that if a write - request has been initiated no read - requests should be latched unless the
  write - response has arrived.
  The contraint is fullilled using the register wr_write_req which holds the current address of
  the line being written to the fabric on a eviction. When such a conflict is detected we store the
  popped request from the data memory subsystem into the rg_read_line_req register so that it can be
  handled once the conflict is done.
  */
  rule rl_handle_dmem_line_read_request(rg_read_line_req matches tagged Invalid );
    Bool perform_req = True;
  	let req <- dmem.send_mem_rd_req.get;
	AXI4_Rd_Addr#(`paddr,`axi4_id_width, 0) dmem_request = AXI4_Rd_Addr {araddr : truncate(req.address), aruser: ?,
      arlen : req.burst_len, arsize : req.burst_size, arburst : 'b10, // arburst : 00 - FIXED 01 - INCR 10 - WRAP
      arid : 0 ,arprot:{1'b0, 1'b0, curr_priv[1]} }; 
    if(wr_write_req matches tagged Valid .waddr) begin
      if((waddr>>(`dwords + `dblocks )) == (req.address>>(`dwords + `dblocks ) ))begin
        perform_req = False;
        rg_read_line_req <= tagged Valid dmem_request;
        `logLevel( core, 1, $format("[%2d]CORE: Delaying Request: ",hartid,fshow(req)))
      end
    end
    if(perform_req)  begin
 	    memory_xactor.i_rd_addr.enq(dmem_request);
      `logLevel( core, 1, $format("[%2d]CORE : DMEM Line Requesting ",hartid, fshow(dmem_request)))
    end
	endrule:rl_handle_dmem_line_read_request

  /*doc:rule: This rule will fire when a pending read operation is present due to a RAW conflict on
   * the line address*/
  rule rl_handle_delayed_read(rg_read_line_req matches tagged Valid .r &&& 
                                  wr_write_req matches tagged Invalid );
	  memory_xactor.i_rd_addr.enq(r);
    `logLevel( core, 1, $format("[%2d]CORE : DMEM Delayed Line Requesting ",hartid, fshow(r)))
    rg_read_line_req <= tagged Invalid;
  endrule:rl_handle_delayed_read

	rule rl_handle_dmem_line_resp(memory_xactor.o_rd_data.first.rid == 0);
    let fab_resp <- pop_o (memory_xactor.o_rd_data);
		let lv_data= fab_resp.rdata;
  	Bool bus_error = !(fab_resp.rresp == AXI4_OKAY); 
    dmem.receive_mem_rd_resp.put(DCache_mem_readresp{data:truncate(lv_data),
                                               last:fab_resp.rlast,
                                               err :bus_error});
    `logLevel( core, 1, $format("[%2d]CORE : DMEM Line Response ",hartid, fshow(fab_resp)))
  endrule:rl_handle_dmem_line_resp

  /*doc:rule: This rule is fired when the data memory subsytem is requesting to write an entire line
   * back to memory. This rule will only fire if both the write address channel and the write data
  * channel are capable of taking in new transactions. In this rule we will enqueue the first beat
  * of line. Once sent, the rg_burst_count count is incremented preventing this rule from firing in
  * the susequent cycles untill all the beats of the line has been delivered.*/
  rule rl_handle_dmem_write_request (rg_burst_count == 0);
    // pop the request from the data cache.
    let req = dmem.send_mem_wr_req;

    // write strobe will always be all-ones.
	  Bit#(TDiv#(`buswidth, 8)) write_strobe = '1;

  	// increment burst count to indicate one beat has been sent.
      rg_burst_count <= rg_burst_count + 1;

      AXI4_Wr_Addr#(`paddr,`axi4_id_width, 0) aw = AXI4_Wr_Addr {awaddr : truncate(req.address), awuser : 0,
      awlen : req.burst_len, awsize : zeroExtend(req.burst_size), awburst : 'b01,
      awid : 0, awprot:{1'b0, 1'b0, curr_priv[1]} }; // arburst : 00 - FIXED 01 - INCR 10 - WRAP

	  let w  = AXI4_Wr_Data {wdata : truncate(req.data), wstrb : write_strobe,
                           wlast : req.burst_len == 0, 
                           wid : 0};
    memory_xactor.i_wr_addr.enq(aw);
	  memory_xactor.i_wr_data.enq(w);
    `logLevel( core, 1, $format("[%2d]CORE : DMEM Line Write Addr : Request ",hartid, fshow(aw)))
    if(req.burst_len != 0 )
      wr_write_req <= tagged Valid req.address;
  endrule:rl_handle_dmem_write_request

  /*doc:rule: This rule sends the burst beats of the line write operation. On each iteration the
  * line is read from the eviction fifo of the data memory subystem and shifted by an appropriate
  * amount indicating the beat number. On the last beat, the eviction fifo is dequence and the burst
  * counter is reset to zero. We also invalidate the wr_write_req register on the last beat*/
  rule rl_dmem_burst_write_data(rg_burst_count != 0);
    // last beat is detected if the burst_counter has reached the size of the words in each line -1.
    Bool last = rg_burst_count == fromInteger(((`dblocks * `dwords * 8) / `buswidth)  - 1 );

    // read the eviction fifo
    let req = dmem.send_mem_wr_req;

    // shift line by the relevant the amount
    req.data = req.data >> rg_shift_amount;
	  let w  = AXI4_Wr_Data {wdata : truncate(req.data), wstrb : '1, wlast : last,
                           wid : 0};
    Bit#(TAdd#(TAdd#(TLog#(`dwords), 1), 3)) shift = {`dwords, 3'b0};

    // if last reset all state and exit this loop
    if(last) begin
      rg_burst_count <= 0;
      rg_shift_amount <= `buswidth;
      wr_write_req <= tagged Invalid;
      dmem.deq_mem_wr_req;
    end
    else begin
      // generate the next shift amount and increment rg_burst_count counter.
      rg_shift_amount <= rg_shift_amount + `buswidth;
      rg_burst_count <= rg_burst_count + 1;
    end
	  memory_xactor.i_wr_data.enq(w);
    `logLevel( core, 1, $format("[%2d]CORE : DMEM Write Data: %h rg_burst_count: %d last: %b \
_shift_amount:%d",hartid, req.data, rg_burst_count, last, rg_shift_amount))
  endrule:rl_dmem_burst_write_data

  /*doc:rule: This rule will simply forward the response obtained from the fabric for a previous
   * line write operation to the data memory subsystem*/
  rule handle_dmem_line_write_resp (memory_xactor.o_wr_resp.first.bid == 0);
    let response <- pop_o(memory_xactor.o_wr_resp);
  	let bus_error = !(response.bresp == AXI4_OKAY);
	  dmem.receive_mem_wr_resp.put(bus_error);
    `logLevel( core, 1, $format("[%2d]CORE : DMEM Write Line Response ",hartid, fshow(response)))
  endrule: handle_dmem_line_write_resp

`ifdef itim 
  rule handle_dmem_itim_read_response;
  	let response <- imem.get_mem_read_itim_resp.get;
  	Bool bus_error = response.err;
    dmem.put_nc_read_resp.put(DCache_mem_readresp{data:zeroExtend(response.data),
                                              last:True,
                                              err :bus_error});
    `logLevel( core, 1, $format("[%2d]CORE : DMEM ITIM Response ",hartid, fshow(response)))
  endrule
  rule handle_itim_write_resp;
  	let response <- imem.get_mem_write_itim_resp.get;
  	Bool bus_error = response;
  	riscv.s5_cache.ma_io_response(tagged Valid tuple2(pack(bus_error),?));
    `logLevel( core, 1, $format("[%2d]CORE : ITIM Memory Write Response ",hartid, fshow(response)))
  endrule
`endif
`endif

  mkConnection(imem.ma_curr_priv, curr_priv);
  mkConnection(dmem.ma_curr_priv, curr_priv);

`ifdef supervisor
  // if supervisor is implemented connect the various csrs required by the ptwalk and dtlb modules
  // here
  mkConnection(imem.ma_satp_from_csr,riscv.csrs.mv_csr_satp);
  mkConnection(dmem.ma_satp_from_csr, riscv.csrs.mv_csr_satp);
  mkConnection(dmem.ma_mstatus_from_csr, riscv.csrs.mv_csr_mstatus);
  mkConnection(ptwalk.ma_satp_from_csr,riscv.csrs.mv_csr_satp);
  mkConnection(ptwalk.ma_mstatus_from_csr, riscv.csrs.mv_csr_mstatus);
  `ifndef hypervisor
  mkConnection(ptwalk.ma_curr_priv,curr_priv);
  `endif
  `ifdef hypervisor
    mkConnection(ptwalk.ma_hgatp_from_csr,riscv.csrs.mv_csr_hgatp);
    mkConnection(ptwalk.ma_vsatp_from_csr,riscv.csrs.mv_csr_vsatp);
    mkConnection(ptwalk.ma_hstatus_from_csr, riscv.csrs.mv_csr_hstatus);
    mkConnection(ptwalk.ma_vsstatus_from_csr, riscv.csrs.mv_csr_vsstatus);
    mkConnection(dmem.ma_vsatp_from_csr,riscv.csrs.mv_csr_vsatp);
    mkConnection(dmem.ma_vsstatus_from_csr, riscv.csrs.mv_csr_vsstatus);
    mkConnection(imem.ma_vsatp_from_csr,riscv.csrs.mv_csr_vsatp);
    mkConnection(imem.ma_vs_mode, riscv.csrs.mv_vs_bit);				//vs_bit from from csr_grp1		
  `endif
  /*doc:rule: this rule forwards the tlb miss request from the itlb to the pagetable walk module.
  * This only fires if the page-table walk module is not already handling a miss*/
  rule rl_itlb_req_to_ptwalk(rg_ptw_state == None);
    let req <- imem.get_request_to_ptw.get();
    ptwalk.from_tlb.put(req);
    rg_ptw_state <= IWalk;
  endrule:rl_itlb_req_to_ptwalk

  /*doc:rule: This rule passes the response from the ptwalk-module to the itlb*/
  rule rl_ptwalk_resp_to_itlb(rg_ptw_state == IWalk);
    let resp <- ptwalk.to_tlb.get();
    imem.put_response_frm_ptw.put(resp);
    rg_ptw_state <= None;
  endrule:rl_ptwalk_resp_to_itlb

  /*doc:rule: This rule is used to connect the request from the data tlb to the ptwalk-module. Fires
   * only when the ptwalk is not already processing another tlb miss*/
  rule rl_dtlb_req_to_ptwalk(rg_ptw_state == None);
    let req <- dmem.get_req_to_ptw.get();
    ptwalk.from_tlb.put(req);
    rg_ptw_state <= DWalk;
  endrule:rl_dtlb_req_to_ptwalk

  /*doc:rule: This rule connects the ptwalk-module response to the data tlb*/
  rule rl_ptwalk_resp_to_dtlb(rg_ptw_state == DWalk);
    let resp <- ptwalk.to_tlb.get();
    dmem.put_resp_from_ptw.put(resp);
    rg_ptw_state <= None;
  endrule:rl_ptwalk_resp_to_dtlb

  /*doc:connect: this connects the ptwalk request to the data memory subsystem*/
  let ptwalk_req <- mkConnection(dmem.receive_core_req, ptwalk.request_to_cache);

  /*doc:connect: This connects the data memory response to the ptwalk-module*/
  mkConnection(dmem.get_ptw_resp, ptwalk.response_frm_cache);

  /*doc:connect: when a tlb-miss occurs in the data tlb, we need to park the original request in the
   * ptwalk-module so that it can be replayed again at the end of the walk.*/
  mkConnection(dmem.get_hold_req, ptwalk.hold_req);
`endif
`ifdef perfmonitors
  `ifdef icache
    mkConnection(riscv.perfmonitors.ma_icache_counters,imem.mv_icache_perf_counters);
  `endif
  `ifdef dcache
    mkConnection(riscv.perfmonitors.ma_dcache_counters,dmem.mv_dcache_perf_counters);
  `endif
  `ifdef supervisor
    mkConnection(riscv.perfmonitors.ma_itlb_counters,imem.mv_itlb_perf_counters);
    mkConnection(riscv.perfmonitors.ma_dtlb_counters,dmem.mv_dtlb_perf_counters);
  `endif
`endif   
  interface sb_clint_msip = interface Put
    method Action put(Bit#(1) intrpt);
      riscv.interrupts.ma_clint_msip(intrpt);
    endmethod
  endinterface;
  interface sb_clint_mtip = interface Put
    method Action put(Bit#(1) intrpt);
      riscv.interrupts.ma_clint_mtip(intrpt);
    endmethod
  endinterface;
  interface sb_clint_mtime = interface Put
    method Action put (Bit#(64) c_mtime);
      riscv.interrupts.ma_clint_mtime(c_mtime);
    endmethod
  endinterface;
	method sb_plic_meip  = riscv.interrupts.ma_plic_meip;
`ifdef supervisor
	method sb_plic_seip = riscv.interrupts.ma_plic_seip;
`endif
`ifdef usertraps
	method sb_plic_ueip = riscv.interrupts.ma_plic_ueip;
`endif
	interface master_i = fetch_xactor.axi_side;
	interface master_d = memory_xactor.axi_side;
`ifdef rtldump
  interface commitlog = riscv.commitlog;
  interface sbread = riscv.sbread;
`endif
`ifdef debug
  method ma_debug_interrupt= riscv.ma_debug_interrupt;
  method mv_core_is_reset = riscv.mv_core_is_reset;
  method mv_core_debugenable = riscv.mv_core_debugenable;
  method ma_debugger_available = riscv.ma_debugger_available;
  method mv_stop_timer = riscv.mv_stop_timer;
  method mv_stop_count = riscv.mv_stop_count;
`endif
endmodule : mkccore_axi4
endpackage:ccore
